/*
$\varphi(n)$ for $M_{ZC}=12$
u φ(0),…,φ(11)

*/
module varphi12 (
    input [4:0] i_u,  //! 0,1,...,29      (sequence group)
    input [3:0] i_n,  //! 0,1,...,M_ZC-1 = 11  (index of φ)

    output [PHI_EN_BITS-1:0] o_varphi_n  // 10 11 00 01 ~ -3 -1 1 3 φ(n)
);

  localparam PHI_EN_BITS = 02;  // Varphi encode define
  localparam PHI_EN_NUMS = 12;  // Varphi encode define
  localparam PHI_EN_NEG_3 = 2'b10;  // Varphi encode define
  localparam PHI_EN_NEG_1 = 2'b11;  // Varphi encode define
  localparam PHI_EN_POS_1 = 2'b00;  // Varphi encode define
  localparam PHI_EN_POS_3 = 2'b01;  // Varphi encode define

  // Declaration of the 2D array
  wire [PHI_EN_NUMS * PHI_EN_BITS-1:0] varphi[0:29];

  //     varphi[u]  =  φ(n) n \in {0,1,...,M_ZC-1}
  assign varphi[0]  = {PHI_EN_NEG_3, PHI_EN_POS_1, PHI_EN_NEG_3, PHI_EN_NEG_3, PHI_EN_NEG_3, PHI_EN_POS_3, PHI_EN_NEG_3, PHI_EN_NEG_1, PHI_EN_POS_1, PHI_EN_POS_1, PHI_EN_POS_1, PHI_EN_NEG_3};
  assign varphi[1]  = {PHI_EN_NEG_3, PHI_EN_POS_3, PHI_EN_POS_1, PHI_EN_NEG_3, PHI_EN_POS_1, PHI_EN_POS_3, PHI_EN_NEG_1, PHI_EN_NEG_1, PHI_EN_POS_1, PHI_EN_POS_3, PHI_EN_POS_3, PHI_EN_POS_3};
  assign varphi[2]  = {PHI_EN_NEG_3, PHI_EN_POS_3, PHI_EN_POS_3, PHI_EN_POS_1, PHI_EN_NEG_3, PHI_EN_POS_3, PHI_EN_NEG_1, PHI_EN_POS_1, PHI_EN_POS_3, PHI_EN_NEG_3, PHI_EN_POS_3, PHI_EN_NEG_3};
  assign varphi[3]  = {PHI_EN_NEG_3, PHI_EN_NEG_3, PHI_EN_NEG_1, PHI_EN_POS_3, PHI_EN_POS_3, PHI_EN_POS_3, PHI_EN_NEG_3, PHI_EN_POS_3, PHI_EN_NEG_3, PHI_EN_POS_1, PHI_EN_NEG_1, PHI_EN_NEG_3};
  assign varphi[4]  = {PHI_EN_NEG_3, PHI_EN_NEG_1, PHI_EN_NEG_1, PHI_EN_POS_1, PHI_EN_POS_3, PHI_EN_POS_1, PHI_EN_POS_1, PHI_EN_NEG_1, PHI_EN_POS_1, PHI_EN_NEG_1, PHI_EN_NEG_3, PHI_EN_POS_1};
  assign varphi[5]  = {PHI_EN_NEG_3, PHI_EN_NEG_3, PHI_EN_POS_3, PHI_EN_POS_1, PHI_EN_NEG_3, PHI_EN_NEG_3, PHI_EN_NEG_3, PHI_EN_NEG_1, PHI_EN_POS_3, PHI_EN_NEG_1, PHI_EN_POS_1, PHI_EN_POS_3};
  assign varphi[6]  = {PHI_EN_POS_1, PHI_EN_NEG_1, PHI_EN_POS_3, PHI_EN_NEG_1, PHI_EN_NEG_1, PHI_EN_NEG_1, PHI_EN_NEG_3, PHI_EN_NEG_1, PHI_EN_POS_1, PHI_EN_POS_1, PHI_EN_POS_1, PHI_EN_NEG_3};
  assign varphi[7]  = {PHI_EN_NEG_1, PHI_EN_NEG_3, PHI_EN_POS_3, PHI_EN_NEG_1, PHI_EN_NEG_3, PHI_EN_NEG_3, PHI_EN_NEG_3, PHI_EN_NEG_1, PHI_EN_POS_1, PHI_EN_NEG_1, PHI_EN_POS_1, PHI_EN_NEG_3};
  assign varphi[8]  = {PHI_EN_NEG_3, PHI_EN_NEG_1, PHI_EN_POS_3, PHI_EN_POS_1, PHI_EN_NEG_3, PHI_EN_NEG_1, PHI_EN_NEG_3, PHI_EN_POS_3, PHI_EN_POS_1, PHI_EN_POS_3, PHI_EN_POS_3, PHI_EN_POS_1};
  assign varphi[9]  = {PHI_EN_NEG_3, PHI_EN_NEG_1, PHI_EN_NEG_1, PHI_EN_NEG_3, PHI_EN_NEG_3, PHI_EN_NEG_1, PHI_EN_NEG_3, PHI_EN_POS_3, PHI_EN_POS_1, PHI_EN_POS_3, PHI_EN_NEG_1, PHI_EN_NEG_3};
  assign varphi[10] = {PHI_EN_NEG_3, PHI_EN_POS_3, PHI_EN_NEG_3, PHI_EN_POS_3, PHI_EN_POS_3, PHI_EN_NEG_3, PHI_EN_NEG_1, PHI_EN_NEG_1, PHI_EN_POS_3, PHI_EN_POS_3, PHI_EN_POS_1, PHI_EN_NEG_3};
  assign varphi[11] = {PHI_EN_NEG_3, PHI_EN_NEG_1, PHI_EN_NEG_3, PHI_EN_NEG_1, PHI_EN_NEG_1, PHI_EN_NEG_3, PHI_EN_POS_3, PHI_EN_POS_3, PHI_EN_NEG_1, PHI_EN_NEG_1, PHI_EN_POS_1, PHI_EN_NEG_3};
  assign varphi[12] = {PHI_EN_NEG_3, PHI_EN_NEG_1, PHI_EN_POS_3, PHI_EN_NEG_3, PHI_EN_NEG_3, PHI_EN_NEG_1, PHI_EN_NEG_3, PHI_EN_POS_1, PHI_EN_NEG_1, PHI_EN_NEG_3, PHI_EN_POS_3, PHI_EN_POS_3};
  assign varphi[13] = {PHI_EN_NEG_3, PHI_EN_POS_1, PHI_EN_NEG_1, PHI_EN_NEG_1, PHI_EN_POS_3, PHI_EN_POS_3, PHI_EN_NEG_3, PHI_EN_NEG_1, PHI_EN_NEG_1, PHI_EN_NEG_3, PHI_EN_NEG_1, PHI_EN_NEG_3};
  assign varphi[14] = {PHI_EN_POS_1, PHI_EN_POS_3, PHI_EN_NEG_3, PHI_EN_POS_1, PHI_EN_POS_3, PHI_EN_POS_3, PHI_EN_POS_3, PHI_EN_POS_1, PHI_EN_NEG_1, PHI_EN_POS_1, PHI_EN_NEG_1, PHI_EN_POS_3};
  assign varphi[15] = {PHI_EN_NEG_3, PHI_EN_POS_1, PHI_EN_POS_3, PHI_EN_NEG_1, PHI_EN_NEG_1, PHI_EN_NEG_3, PHI_EN_NEG_3, PHI_EN_NEG_1, PHI_EN_NEG_1, PHI_EN_POS_3, PHI_EN_POS_1, PHI_EN_NEG_3};
  assign varphi[16] = {PHI_EN_NEG_1, PHI_EN_NEG_1, PHI_EN_NEG_1, PHI_EN_NEG_1, PHI_EN_POS_1, PHI_EN_NEG_3, PHI_EN_NEG_1, PHI_EN_POS_3, PHI_EN_POS_3, PHI_EN_NEG_1, PHI_EN_NEG_3, PHI_EN_POS_1};
  assign varphi[17] = {PHI_EN_NEG_1, PHI_EN_POS_1, PHI_EN_POS_1, PHI_EN_NEG_1, PHI_EN_POS_1, PHI_EN_POS_3, PHI_EN_POS_3, PHI_EN_NEG_1, PHI_EN_NEG_1, PHI_EN_NEG_3, PHI_EN_POS_1, PHI_EN_NEG_3};
  assign varphi[18] = {PHI_EN_NEG_3, PHI_EN_POS_1, PHI_EN_POS_3, PHI_EN_POS_3, PHI_EN_NEG_1, PHI_EN_NEG_1, PHI_EN_NEG_3, PHI_EN_POS_3, PHI_EN_POS_3, PHI_EN_NEG_3, PHI_EN_POS_3, PHI_EN_NEG_3};
  assign varphi[19] = {PHI_EN_NEG_3, PHI_EN_NEG_3, PHI_EN_POS_3, PHI_EN_NEG_3, PHI_EN_NEG_1, PHI_EN_POS_3, PHI_EN_POS_3, PHI_EN_POS_3, PHI_EN_NEG_1, PHI_EN_NEG_3, PHI_EN_POS_1, PHI_EN_NEG_3};
  assign varphi[20] = {PHI_EN_POS_3, PHI_EN_POS_1, PHI_EN_POS_3, PHI_EN_POS_1, PHI_EN_POS_3, PHI_EN_NEG_3, PHI_EN_NEG_1, PHI_EN_POS_1, PHI_EN_POS_3, PHI_EN_POS_1, PHI_EN_NEG_1, PHI_EN_NEG_3};
  assign varphi[21] = {PHI_EN_NEG_3, PHI_EN_POS_3, PHI_EN_POS_1, PHI_EN_POS_3, PHI_EN_NEG_3, PHI_EN_POS_1, PHI_EN_POS_1, PHI_EN_POS_1, PHI_EN_POS_1, PHI_EN_POS_3, PHI_EN_NEG_3, PHI_EN_POS_3};
  assign varphi[22] = {PHI_EN_NEG_3, PHI_EN_POS_3, PHI_EN_POS_3, PHI_EN_POS_3, PHI_EN_NEG_1, PHI_EN_NEG_3, PHI_EN_NEG_3, PHI_EN_NEG_1, PHI_EN_NEG_3, PHI_EN_POS_1, PHI_EN_POS_3, PHI_EN_NEG_3};
  assign varphi[23] = {PHI_EN_POS_3, PHI_EN_NEG_1, PHI_EN_NEG_3, PHI_EN_POS_3, PHI_EN_NEG_3, PHI_EN_NEG_1, PHI_EN_POS_3, PHI_EN_POS_3, PHI_EN_POS_3, PHI_EN_NEG_3, PHI_EN_NEG_1, PHI_EN_NEG_3};
  assign varphi[24] = {PHI_EN_NEG_3, PHI_EN_NEG_1, PHI_EN_POS_1, PHI_EN_NEG_3, PHI_EN_POS_1, PHI_EN_POS_3, PHI_EN_POS_3, PHI_EN_POS_3, PHI_EN_NEG_1, PHI_EN_NEG_3, PHI_EN_POS_3, PHI_EN_POS_3};
  assign varphi[25] = {PHI_EN_NEG_3, PHI_EN_POS_3, PHI_EN_POS_1, PHI_EN_NEG_1, PHI_EN_POS_3, PHI_EN_POS_3, PHI_EN_NEG_3, PHI_EN_POS_1, PHI_EN_NEG_1, PHI_EN_POS_1, PHI_EN_NEG_1, PHI_EN_POS_1};
  assign varphi[26] = {PHI_EN_NEG_1, PHI_EN_POS_1, PHI_EN_POS_3, PHI_EN_NEG_3, PHI_EN_POS_1, PHI_EN_NEG_1, PHI_EN_POS_1, PHI_EN_NEG_1, PHI_EN_NEG_1, PHI_EN_NEG_3, PHI_EN_POS_1, PHI_EN_NEG_1};
  assign varphi[27] = {PHI_EN_NEG_3, PHI_EN_NEG_3, PHI_EN_POS_3, PHI_EN_POS_3, PHI_EN_POS_3, PHI_EN_NEG_3, PHI_EN_NEG_1, PHI_EN_POS_1, PHI_EN_NEG_3, PHI_EN_POS_3, PHI_EN_POS_1, PHI_EN_NEG_3};
  assign varphi[28] = {PHI_EN_POS_1, PHI_EN_NEG_1, PHI_EN_POS_3, PHI_EN_POS_1, PHI_EN_POS_1, PHI_EN_NEG_1, PHI_EN_NEG_1, PHI_EN_NEG_1, PHI_EN_POS_1, PHI_EN_POS_3, PHI_EN_NEG_3, PHI_EN_POS_1};
  assign varphi[29] = {PHI_EN_NEG_3, PHI_EN_POS_3, PHI_EN_NEG_3, PHI_EN_POS_3, PHI_EN_NEG_3, PHI_EN_NEG_3, PHI_EN_POS_3, PHI_EN_NEG_1, PHI_EN_NEG_1, PHI_EN_POS_1, PHI_EN_POS_3, PHI_EN_NEG_3};


  // wire [31:0] test = {i_n, {(`PHI_EN_BITS - 1){1'b0}}};
  wire [PHI_EN_NUMS*PHI_EN_BITS-1:0] varphi_shift = varphi[i_u] << {i_n, {(PHI_EN_BITS - 1) {1'b0}}};  // shift by number of varphi encode bits

  assign o_varphi_n = varphi_shift[PHI_EN_NUMS*PHI_EN_BITS-1:(PHI_EN_NUMS-1)*PHI_EN_BITS];

endmodule
