/*
    Point  1: Real = 0111111111111111 (1.0000), Imaginary = 0000000000000000 (0.0000)
    Point  2: Real = 0111111111101110 (0.9995), Imaginary = 0000010000110000 (0.0327)
    Point  3: Real = 0111111110111010 (0.9979), Imaginary = 0000100001011111 (0.0654)
    Point  4: Real = 0111111101100010 (0.9952), Imaginary = 0000110010001100 (0.0980)
    Point  5: Real = 0111111011101000 (0.9914), Imaginary = 0001000010110101 (0.1305)
    Point  6: Real = 0111111001001010 (0.9866), Imaginary = 0001010011011010 (0.1629)
    Point  7: Real = 0111110110001010 (0.9808), Imaginary = 0001100011111001 (0.1951)
    Point  8: Real = 0111110010101000 (0.9739), Imaginary = 0001110100010001 (0.2271)
    Point  9: Real = 0111101110100011 (0.9659), Imaginary = 0010000100100001 (0.2588)
    Point 10: Real = 0111101001111101 (0.9569), Imaginary = 0010010100101000 (0.2903)
    Point 11: Real = 0111100100110101 (0.9469), Imaginary = 0010100100100101 (0.3214)
    Point 12: Real = 0111011111001100 (0.9359), Imaginary = 0010110100010111 (0.3523)
    Point 13: Real = 0111011001000010 (0.9239), Imaginary = 0011000011111100 (0.3827)
    Point 14: Real = 0111010010010111 (0.9109), Imaginary = 0011010011010100 (0.4127)
    Point 15: Real = 0111001011001101 (0.8969), Imaginary = 0011100010011101 (0.4423)
    Point 16: Real = 0111000011100011 (0.8819), Imaginary = 0011110001010111 (0.4714)
    Point 17: Real = 0110111011011010 (0.8660), Imaginary = 0100000000000000 (0.5000)
    Point 18: Real = 0110110010110011 (0.8492), Imaginary = 0100001110011000 (0.5281)
    Point 19: Real = 0110101001101110 (0.8315), Imaginary = 0100011100011101 (0.5556)
    Point 20: Real = 0110100000001011 (0.8128), Imaginary = 0100101010001111 (0.5825)
    Point 21: Real = 0110010110001101 (0.7934), Imaginary = 0100110111101100 (0.6088)
    Point 22: Real = 0110001011110010 (0.7730), Imaginary = 0101000100110100 (0.6344)
    Point 23: Real = 0110000000111100 (0.7518), Imaginary = 0101010001100101 (0.6593)
    Point 24: Real = 0101110101101100 (0.7299), Imaginary = 0101011110000000 (0.6836)
    Point 25: Real = 0101101010000010 (0.7071), Imaginary = 0101101010000010 (0.7071)
    Point 26: Real = 0101011110000000 (0.6836), Imaginary = 0101110101101100 (0.7299)
    Point 27: Real = 0101010001100101 (0.6593), Imaginary = 0110000000111100 (0.7518)
    Point 28: Real = 0101000100110100 (0.6344), Imaginary = 0110001011110010 (0.7730)
    Point 29: Real = 0100110111101100 (0.6088), Imaginary = 0110010110001101 (0.7934)
    Point 30: Real = 0100101010001111 (0.5825), Imaginary = 0110100000001011 (0.8128)
    Point 31: Real = 0100011100011101 (0.5556), Imaginary = 0110101001101110 (0.8315)
    Point 32: Real = 0100001110011000 (0.5281), Imaginary = 0110110010110011 (0.8492)
    Point 33: Real = 0100000000000000 (0.5000), Imaginary = 0110111011011010 (0.8660)
    Point 34: Real = 0011110001010111 (0.4714), Imaginary = 0111000011100011 (0.8819)
    Point 35: Real = 0011100010011101 (0.4423), Imaginary = 0111001011001101 (0.8969)
    Point 36: Real = 0011010011010100 (0.4127), Imaginary = 0111010010010111 (0.9109)
    Point 37: Real = 0011000011111100 (0.3827), Imaginary = 0111011001000010 (0.9239)
    Point 38: Real = 0010110100010111 (0.3523), Imaginary = 0111011111001100 (0.9359)
    Point 39: Real = 0010100100100101 (0.3214), Imaginary = 0111100100110101 (0.9469)
    Point 40: Real = 0010010100101000 (0.2903), Imaginary = 0111101001111101 (0.9569)
    Point 41: Real = 0010000100100001 (0.2588), Imaginary = 0111101110100011 (0.9659)
    Point 42: Real = 0001110100010001 (0.2271), Imaginary = 0111110010101000 (0.9739)
    Point 43: Real = 0001100011111001 (0.1951), Imaginary = 0111110110001010 (0.9808)
    Point 44: Real = 0001010011011010 (0.1629), Imaginary = 0111111001001010 (0.9866)
    Point 45: Real = 0001000010110101 (0.1305), Imaginary = 0111111011101000 (0.9914)
    Point 46: Real = 0000110010001100 (0.0980), Imaginary = 0111111101100010 (0.9952)
    Point 47: Real = 0000100001011111 (0.0654), Imaginary = 0111111110111010 (0.9979)
    Point 48: Real = 0000010000110000 (0.0327), Imaginary = 0111111111101110 (0.9995)
    Point 49: Real = 0000000000000000 (0.0000), Imaginary = 0111111111111111 (1.0000)
    Point 50: Real = 1111101111010000 (-0.0327), Imaginary = 0111111111101110 (0.9995)
    Point 51: Real = 1111011110100001 (-0.0654), Imaginary = 0111111110111010 (0.9979)
    Point 52: Real = 1111001101110100 (-0.0980), Imaginary = 0111111101100010 (0.9952)
    Point 53: Real = 1110111101001011 (-0.1305), Imaginary = 0111111011101000 (0.9914)
    Point 54: Real = 1110101100100110 (-0.1629), Imaginary = 0111111001001010 (0.9866)
    Point 55: Real = 1110011100000111 (-0.1951), Imaginary = 0111110110001010 (0.9808)
    Point 56: Real = 1110001011101111 (-0.2271), Imaginary = 0111110010101000 (0.9739)
    Point 57: Real = 1101111011011111 (-0.2588), Imaginary = 0111101110100011 (0.9659)
    Point 58: Real = 1101101011011000 (-0.2903), Imaginary = 0111101001111101 (0.9569)
    Point 59: Real = 1101011011011011 (-0.3214), Imaginary = 0111100100110101 (0.9469)
    Point 60: Real = 1101001011101001 (-0.3523), Imaginary = 0111011111001100 (0.9359)
    Point 61: Real = 1100111100000100 (-0.3827), Imaginary = 0111011001000010 (0.9239)
    Point 62: Real = 1100101100101100 (-0.4127), Imaginary = 0111010010010111 (0.9109)
    Point 63: Real = 1100011101100011 (-0.4423), Imaginary = 0111001011001101 (0.8969)
    Point 64: Real = 1100001110101001 (-0.4714), Imaginary = 0111000011100011 (0.8819)
    Point 65: Real = 1100000000000000 (-0.5000), Imaginary = 0110111011011010 (0.8660)
    Point 66: Real = 1011110001101000 (-0.5281), Imaginary = 0110110010110011 (0.8492)
    Point 67: Real = 1011100011100011 (-0.5556), Imaginary = 0110101001101110 (0.8315)
    Point 68: Real = 1011010101110001 (-0.5825), Imaginary = 0110100000001011 (0.8128)
    Point 69: Real = 1011001000010100 (-0.6088), Imaginary = 0110010110001101 (0.7934)
    Point 70: Real = 1010111011001100 (-0.6344), Imaginary = 0110001011110010 (0.7730)
    Point 71: Real = 1010101110011011 (-0.6593), Imaginary = 0110000000111100 (0.7518)
    Point 72: Real = 1010100010000000 (-0.6836), Imaginary = 0101110101101100 (0.7299)
    Point 73: Real = 1010010101111110 (-0.7071), Imaginary = 0101101010000010 (0.7071)
    Point 74: Real = 1010001010010100 (-0.7299), Imaginary = 0101011110000000 (0.6836)
    Point 75: Real = 1001111111000100 (-0.7518), Imaginary = 0101010001100101 (0.6593)
    Point 76: Real = 1001110100001110 (-0.7730), Imaginary = 0101000100110100 (0.6344)
    Point 77: Real = 1001101001110011 (-0.7934), Imaginary = 0100110111101100 (0.6088)
    Point 78: Real = 1001011111110101 (-0.8128), Imaginary = 0100101010001111 (0.5825)
    Point 79: Real = 1001010110010010 (-0.8315), Imaginary = 0100011100011101 (0.5556)
    Point 80: Real = 1001001101001101 (-0.8492), Imaginary = 0100001110011000 (0.5281)
    Point 81: Real = 1001000100100110 (-0.8660), Imaginary = 0100000000000000 (0.5000)
    Point 82: Real = 1000111100011101 (-0.8819), Imaginary = 0011110001010111 (0.4714)
    Point 83: Real = 1000110100110011 (-0.8969), Imaginary = 0011100010011101 (0.4423)
    Point 84: Real = 1000101101101001 (-0.9109), Imaginary = 0011010011010100 (0.4127)
    Point 85: Real = 1000100110111110 (-0.9239), Imaginary = 0011000011111100 (0.3827)
    Point 86: Real = 1000100000110100 (-0.9359), Imaginary = 0010110100010111 (0.3523)
    Point 87: Real = 1000011011001011 (-0.9469), Imaginary = 0010100100100101 (0.3214)
    Point 88: Real = 1000010110000011 (-0.9569), Imaginary = 0010010100101000 (0.2903)
    Point 89: Real = 1000010001011101 (-0.9659), Imaginary = 0010000100100001 (0.2588)
    Point 90: Real = 1000001101011000 (-0.9739), Imaginary = 0001110100010001 (0.2271)
    Point 91: Real = 1000001001110110 (-0.9808), Imaginary = 0001100011111001 (0.1951)
    Point 92: Real = 1000000110110110 (-0.9866), Imaginary = 0001010011011010 (0.1629)
    Point 93: Real = 1000000100011000 (-0.9914), Imaginary = 0001000010110101 (0.1305)
    Point 94: Real = 1000000010011110 (-0.9952), Imaginary = 0000110010001100 (0.0980)
    Point 95: Real = 1000000001000110 (-0.9979), Imaginary = 0000100001011111 (0.0654)
    Point 96: Real = 1000000000010010 (-0.9995), Imaginary = 0000010000110000 (0.0327)
    Point 97: Real = 1000000000000000 (-1.0000), Imaginary = 0000000000000000 (0.0000)
    Point 98: Real = 1000000000010010 (-0.9995), Imaginary = 1111101111010000 (-0.0327)
    Point 99: Real = 1000000001000110 (-0.9979), Imaginary = 1111011110100001 (-0.0654)
    Point 100: Real = 1000000010011110 (-0.9952), Imaginary = 1111001101110100 (-0.0980)
    Point 101: Real = 1000000100011000 (-0.9914), Imaginary = 1110111101001011 (-0.1305)
    Point 102: Real = 1000000110110110 (-0.9866), Imaginary = 1110101100100110 (-0.1629)
    Point 103: Real = 1000001001110110 (-0.9808), Imaginary = 1110011100000111 (-0.1951)
    Point 104: Real = 1000001101011000 (-0.9739), Imaginary = 1110001011101111 (-0.2271)
    Point 105: Real = 1000010001011101 (-0.9659), Imaginary = 1101111011011111 (-0.2588)
    Point 106: Real = 1000010110000011 (-0.9569), Imaginary = 1101101011011000 (-0.2903)
    Point 107: Real = 1000011011001011 (-0.9469), Imaginary = 1101011011011011 (-0.3214)
    Point 108: Real = 1000100000110100 (-0.9359), Imaginary = 1101001011101001 (-0.3523)
    Point 109: Real = 1000100110111110 (-0.9239), Imaginary = 1100111100000100 (-0.3827)
    Point 110: Real = 1000101101101001 (-0.9109), Imaginary = 1100101100101100 (-0.4127)
    Point 111: Real = 1000110100110011 (-0.8969), Imaginary = 1100011101100011 (-0.4423)
    Point 112: Real = 1000111100011101 (-0.8819), Imaginary = 1100001110101001 (-0.4714)
    Point 113: Real = 1001000100100110 (-0.8660), Imaginary = 1100000000000000 (-0.5000)
    Point 114: Real = 1001001101001101 (-0.8492), Imaginary = 1011110001101000 (-0.5281)
    Point 115: Real = 1001010110010010 (-0.8315), Imaginary = 1011100011100011 (-0.5556)
    Point 116: Real = 1001011111110101 (-0.8128), Imaginary = 1011010101110001 (-0.5825)
    Point 117: Real = 1001101001110011 (-0.7934), Imaginary = 1011001000010100 (-0.6088)
    Point 118: Real = 1001110100001110 (-0.7730), Imaginary = 1010111011001100 (-0.6344)
    Point 119: Real = 1001111111000100 (-0.7518), Imaginary = 1010101110011011 (-0.6593)
    Point 120: Real = 1010001010010100 (-0.7299), Imaginary = 1010100010000000 (-0.6836)
    Point 121: Real = 1010010101111110 (-0.7071), Imaginary = 1010010101111110 (-0.7071)
    Point 122: Real = 1010100010000000 (-0.6836), Imaginary = 1010001010010100 (-0.7299)
    Point 123: Real = 1010101110011011 (-0.6593), Imaginary = 1001111111000100 (-0.7518)
    Point 124: Real = 1010111011001100 (-0.6344), Imaginary = 1001110100001110 (-0.7730)
    Point 125: Real = 1011001000010100 (-0.6088), Imaginary = 1001101001110011 (-0.7934)
    Point 126: Real = 1011010101110001 (-0.5825), Imaginary = 1001011111110101 (-0.8128)
    Point 127: Real = 1011100011100011 (-0.5556), Imaginary = 1001010110010010 (-0.8315)
    Point 128: Real = 1011110001101000 (-0.5281), Imaginary = 1001001101001101 (-0.8492)
    Point 129: Real = 1100000000000000 (-0.5000), Imaginary = 1001000100100110 (-0.8660)
    Point 130: Real = 1100001110101001 (-0.4714), Imaginary = 1000111100011101 (-0.8819)
    Point 131: Real = 1100011101100011 (-0.4423), Imaginary = 1000110100110011 (-0.8969)
    Point 132: Real = 1100101100101100 (-0.4127), Imaginary = 1000101101101001 (-0.9109)
    Point 133: Real = 1100111100000100 (-0.3827), Imaginary = 1000100110111110 (-0.9239)
    Point 134: Real = 1101001011101001 (-0.3523), Imaginary = 1000100000110100 (-0.9359)
    Point 135: Real = 1101011011011011 (-0.3214), Imaginary = 1000011011001011 (-0.9469)
    Point 136: Real = 1101101011011000 (-0.2903), Imaginary = 1000010110000011 (-0.9569)
    Point 137: Real = 1101111011011111 (-0.2588), Imaginary = 1000010001011101 (-0.9659)
    Point 138: Real = 1110001011101111 (-0.2271), Imaginary = 1000001101011000 (-0.9739)
    Point 139: Real = 1110011100000111 (-0.1951), Imaginary = 1000001001110110 (-0.9808)
    Point 140: Real = 1110101100100110 (-0.1629), Imaginary = 1000000110110110 (-0.9866)
    Point 141: Real = 1110111101001011 (-0.1305), Imaginary = 1000000100011000 (-0.9914)
    Point 142: Real = 1111001101110100 (-0.0980), Imaginary = 1000000010011110 (-0.9952)
    Point 143: Real = 1111011110100001 (-0.0654), Imaginary = 1000000001000110 (-0.9979)
    Point 144: Real = 1111101111010000 (-0.0327), Imaginary = 1000000000010010 (-0.9995)
    Point 145: Real = 0000000000000000 (-0.0000), Imaginary = 1000000000000000 (-1.0000)
    Point 146: Real = 0000010000110000 (0.0327), Imaginary = 1000000000010010 (-0.9995)
    Point 147: Real = 0000100001011111 (0.0654), Imaginary = 1000000001000110 (-0.9979)
    Point 148: Real = 0000110010001100 (0.0980), Imaginary = 1000000010011110 (-0.9952)
    Point 149: Real = 0001000010110101 (0.1305), Imaginary = 1000000100011000 (-0.9914)
    Point 150: Real = 0001010011011010 (0.1629), Imaginary = 1000000110110110 (-0.9866)
    Point 151: Real = 0001100011111001 (0.1951), Imaginary = 1000001001110110 (-0.9808)
    Point 152: Real = 0001110100010001 (0.2271), Imaginary = 1000001101011000 (-0.9739)
    Point 153: Real = 0010000100100001 (0.2588), Imaginary = 1000010001011101 (-0.9659)
    Point 154: Real = 0010010100101000 (0.2903), Imaginary = 1000010110000011 (-0.9569)
    Point 155: Real = 0010100100100101 (0.3214), Imaginary = 1000011011001011 (-0.9469)
    Point 156: Real = 0010110100010111 (0.3523), Imaginary = 1000100000110100 (-0.9359)
    Point 157: Real = 0011000011111100 (0.3827), Imaginary = 1000100110111110 (-0.9239)
    Point 158: Real = 0011010011010100 (0.4127), Imaginary = 1000101101101001 (-0.9109)
    Point 159: Real = 0011100010011101 (0.4423), Imaginary = 1000110100110011 (-0.8969)
    Point 160: Real = 0011110001010111 (0.4714), Imaginary = 1000111100011101 (-0.8819)
    Point 161: Real = 0100000000000000 (0.5000), Imaginary = 1001000100100110 (-0.8660)
    Point 162: Real = 0100001110011000 (0.5281), Imaginary = 1001001101001101 (-0.8492)
    Point 163: Real = 0100011100011101 (0.5556), Imaginary = 1001010110010010 (-0.8315)
    Point 164: Real = 0100101010001111 (0.5825), Imaginary = 1001011111110101 (-0.8128)
    Point 165: Real = 0100110111101100 (0.6088), Imaginary = 1001101001110011 (-0.7934)
    Point 166: Real = 0101000100110100 (0.6344), Imaginary = 1001110100001110 (-0.7730)
    Point 167: Real = 0101010001100101 (0.6593), Imaginary = 1001111111000100 (-0.7518)
    Point 168: Real = 0101011110000000 (0.6836), Imaginary = 1010001010010100 (-0.7299)
    Point 169: Real = 0101101010000010 (0.7071), Imaginary = 1010010101111110 (-0.7071)
    Point 170: Real = 0101110101101100 (0.7299), Imaginary = 1010100010000000 (-0.6836)
    Point 171: Real = 0110000000111100 (0.7518), Imaginary = 1010101110011011 (-0.6593)
    Point 172: Real = 0110001011110010 (0.7730), Imaginary = 1010111011001100 (-0.6344)
    Point 173: Real = 0110010110001101 (0.7934), Imaginary = 1011001000010100 (-0.6088)
    Point 174: Real = 0110100000001011 (0.8128), Imaginary = 1011010101110001 (-0.5825)
    Point 175: Real = 0110101001101110 (0.8315), Imaginary = 1011100011100011 (-0.5556)
    Point 176: Real = 0110110010110011 (0.8492), Imaginary = 1011110001101000 (-0.5281)
    Point 177: Real = 0110111011011010 (0.8660), Imaginary = 1100000000000000 (-0.5000)
    Point 178: Real = 0111000011100011 (0.8819), Imaginary = 1100001110101001 (-0.4714)
    Point 179: Real = 0111001011001101 (0.8969), Imaginary = 1100011101100011 (-0.4423)
    Point 180: Real = 0111010010010111 (0.9109), Imaginary = 1100101100101100 (-0.4127)
    Point 181: Real = 0111011001000010 (0.9239), Imaginary = 1100111100000100 (-0.3827)
    Point 182: Real = 0111011111001100 (0.9359), Imaginary = 1101001011101001 (-0.3523)
    Point 183: Real = 0111100100110101 (0.9469), Imaginary = 1101011011011011 (-0.3214)
    Point 184: Real = 0111101001111101 (0.9569), Imaginary = 1101101011011000 (-0.2903)
    Point 185: Real = 0111101110100011 (0.9659), Imaginary = 1101111011011111 (-0.2588)
    Point 186: Real = 0111110010101000 (0.9739), Imaginary = 1110001011101111 (-0.2271)
    Point 187: Real = 0111110110001010 (0.9808), Imaginary = 1110011100000111 (-0.1951)
    Point 188: Real = 0111111001001010 (0.9866), Imaginary = 1110101100100110 (-0.1629)
    Point 189: Real = 0111111011101000 (0.9914), Imaginary = 1110111101001011 (-0.1305)
    Point 190: Real = 0111111101100010 (0.9952), Imaginary = 1111001101110100 (-0.0980)
    Point 191: Real = 0111111110111010 (0.9979), Imaginary = 1111011110100001 (-0.0654)
    Point 192: Real = 0111111111101110 (0.9995), Imaginary = 1111101111010000 (-0.0327)
*/

module cyc_192 (
    input [7:0] i_point_index,  //! i_point_index/24 of a cycle (0-191)

    output signed [15:0] o_point_re,  //! Coresponding complex point's real value (sfix16)
    output signed [15:0] o_point_im   //! Coresponding complex point's imaginary value (sfix16)
);

  wire signed [15:0] point_im[0:191];
  wire signed [15:0] point_re[0:191];

  assign o_point_re = point_re[i_point_index];
  assign o_point_im = point_im[i_point_index];

  assign point_re[000] = 'b0111111111111111;  // (1.0000)
  assign point_re[001] = 'b0111111111101110;  // (0.9995)
  assign point_re[002] = 'b0111111110111010;  // (0.9979)
  assign point_re[003] = 'b0111111101100010;  // (0.9952)
  assign point_re[004] = 'b0111111011101000;  // (0.9914)
  assign point_re[005] = 'b0111111001001010;  // (0.9866)
  assign point_re[006] = 'b0111110110001010;  // (0.9808)
  assign point_re[007] = 'b0111110010101000;  // (0.9739)
  assign point_re[008] = 'b0111101110100011;  // (0.9659)
  assign point_re[009] = 'b0111101001111101;  // (0.9569)
  assign point_re[010] = 'b0111100100110101;  // (0.9469)
  assign point_re[011] = 'b0111011111001100;  // (0.9359)
  assign point_re[012] = 'b0111011001000010;  // (0.9239)
  assign point_re[013] = 'b0111010010010111;  // (0.9109)
  assign point_re[014] = 'b0111001011001101;  // (0.8969)
  assign point_re[015] = 'b0111000011100011;  // (0.8819)
  assign point_re[016] = 'b0110111011011010;  // (0.8660)
  assign point_re[017] = 'b0110110010110011;  // (0.8492)
  assign point_re[018] = 'b0110101001101110;  // (0.8315)
  assign point_re[019] = 'b0110100000001011;  // (0.8128)
  assign point_re[020] = 'b0110010110001101;  // (0.7934)
  assign point_re[021] = 'b0110001011110010;  // (0.7730)
  assign point_re[022] = 'b0110000000111100;  // (0.7518)
  assign point_re[023] = 'b0101110101101100;  // (0.7299)
  assign point_re[024] = 'b0101101010000010;  // (0.7071)
  assign point_re[025] = 'b0101011110000000;  // (0.6836)
  assign point_re[026] = 'b0101010001100101;  // (0.6593)
  assign point_re[027] = 'b0101000100110100;  // (0.6344)
  assign point_re[028] = 'b0100110111101100;  // (0.6088)
  assign point_re[029] = 'b0100101010001111;  // (0.5825)
  assign point_re[030] = 'b0100011100011101;  // (0.5556)
  assign point_re[031] = 'b0100001110011000;  // (0.5281)
  assign point_re[032] = 'b0100000000000000;  // (0.5000)
  assign point_re[033] = 'b0011110001010111;  // (0.4714)
  assign point_re[034] = 'b0011100010011101;  // (0.4423)
  assign point_re[035] = 'b0011010011010100;  // (0.4127)
  assign point_re[036] = 'b0011000011111100;  // (0.3827)
  assign point_re[037] = 'b0010110100010111;  // (0.3523)
  assign point_re[038] = 'b0010100100100101;  // (0.3214)
  assign point_re[039] = 'b0010010100101000;  // (0.2903)
  assign point_re[040] = 'b0010000100100001;  // (0.2588)
  assign point_re[041] = 'b0001110100010001;  // (0.2271)
  assign point_re[042] = 'b0001100011111001;  // (0.1951)
  assign point_re[043] = 'b0001010011011010;  // (0.1629)
  assign point_re[044] = 'b0001000010110101;  // (0.1305)
  assign point_re[045] = 'b0000110010001100;  // (0.0980)
  assign point_re[046] = 'b0000100001011111;  // (0.0654)
  assign point_re[047] = 'b0000010000110000;  // (0.0327)
  assign point_re[048] = 'b0000000000000000;  // (0.0000)
  assign point_re[049] = 'b1111101111010000;  // (-0.0327)
  assign point_re[050] = 'b1111011110100001;  // (-0.0654)
  assign point_re[051] = 'b1111001101110100;  // (-0.0980)
  assign point_re[052] = 'b1110111101001011;  // (-0.1305)
  assign point_re[053] = 'b1110101100100110;  // (-0.1629)
  assign point_re[054] = 'b1110011100000111;  // (-0.1951)
  assign point_re[055] = 'b1110001011101111;  // (-0.2271)
  assign point_re[056] = 'b1101111011011111;  // (-0.2588)
  assign point_re[057] = 'b1101101011011000;  // (-0.2903)
  assign point_re[058] = 'b1101011011011011;  // (-0.3214)
  assign point_re[059] = 'b1101001011101001;  // (-0.3523)
  assign point_re[060] = 'b1100111100000100;  // (-0.3827)
  assign point_re[061] = 'b1100101100101100;  // (-0.4127)
  assign point_re[062] = 'b1100011101100011;  // (-0.4423)
  assign point_re[063] = 'b1100001110101001;  // (-0.4714)
  assign point_re[064] = 'b1100000000000000;  // (-0.5000)
  assign point_re[065] = 'b1011110001101000;  // (-0.5281)
  assign point_re[066] = 'b1011100011100011;  // (-0.5556)
  assign point_re[067] = 'b1011010101110001;  // (-0.5825)
  assign point_re[068] = 'b1011001000010100;  // (-0.6088)
  assign point_re[069] = 'b1010111011001100;  // (-0.6344)
  assign point_re[070] = 'b1010101110011011;  // (-0.6593)
  assign point_re[071] = 'b1010100010000000;  // (-0.6836)
  assign point_re[072] = 'b1010010101111110;  // (-0.7071)
  assign point_re[073] = 'b1010001010010100;  // (-0.7299)
  assign point_re[074] = 'b1001111111000100;  // (-0.7518)
  assign point_re[075] = 'b1001110100001110;  // (-0.7730)
  assign point_re[076] = 'b1001101001110011;  // (-0.7934)
  assign point_re[077] = 'b1001011111110101;  // (-0.8128)
  assign point_re[078] = 'b1001010110010010;  // (-0.8315)
  assign point_re[079] = 'b1001001101001101;  // (-0.8492)
  assign point_re[080] = 'b1001000100100110;  // (-0.8660)
  assign point_re[081] = 'b1000111100011101;  // (-0.8819)
  assign point_re[082] = 'b1000110100110011;  // (-0.8969)
  assign point_re[083] = 'b1000101101101001;  // (-0.9109)
  assign point_re[084] = 'b1000100110111110;  // (-0.9239)
  assign point_re[085] = 'b1000100000110100;  // (-0.9359)
  assign point_re[086] = 'b1000011011001011;  // (-0.9469)
  assign point_re[087] = 'b1000010110000011;  // (-0.9569)
  assign point_re[088] = 'b1000010001011101;  // (-0.9659)
  assign point_re[089] = 'b1000001101011000;  // (-0.9739)
  assign point_re[090] = 'b1000001001110110;  // (-0.9808)
  assign point_re[091] = 'b1000000110110110;  // (-0.9866)
  assign point_re[092] = 'b1000000100011000;  // (-0.9914)
  assign point_re[093] = 'b1000000010011110;  // (-0.9952)
  assign point_re[094] = 'b1000000001000110;  // (-0.9979)
  assign point_re[095] = 'b1000000000010010;  // (-0.9995)
  assign point_re[096] = 'b1000000000000000;  // (-1.0000)
  assign point_re[097] = 'b1000000000010010;  // (-0.9995)
  assign point_re[098] = 'b1000000001000110;  // (-0.9979)
  assign point_re[099] = 'b1000000010011110;  // (-0.9952)
  assign point_re[100] = 'b1000000100011000;  // (-0.9914)
  assign point_re[101] = 'b1000000110110110;  // (-0.9866)
  assign point_re[102] = 'b1000001001110110;  // (-0.9808)
  assign point_re[103] = 'b1000001101011000;  // (-0.9739)
  assign point_re[104] = 'b1000010001011101;  // (-0.9659)
  assign point_re[105] = 'b1000010110000011;  // (-0.9569)
  assign point_re[106] = 'b1000011011001011;  // (-0.9469)
  assign point_re[107] = 'b1000100000110100;  // (-0.9359)
  assign point_re[108] = 'b1000100110111110;  // (-0.9239)
  assign point_re[109] = 'b1000101101101001;  // (-0.9109)
  assign point_re[110] = 'b1000110100110011;  // (-0.8969)
  assign point_re[111] = 'b1000111100011101;  // (-0.8819)
  assign point_re[112] = 'b1001000100100110;  // (-0.8660)
  assign point_re[113] = 'b1001001101001101;  // (-0.8492)
  assign point_re[114] = 'b1001010110010010;  // (-0.8315)
  assign point_re[115] = 'b1001011111110101;  // (-0.8128)
  assign point_re[116] = 'b1001101001110011;  // (-0.7934)
  assign point_re[117] = 'b1001110100001110;  // (-0.7730)
  assign point_re[118] = 'b1001111111000100;  // (-0.7518)
  assign point_re[119] = 'b1010001010010100;  // (-0.7299)
  assign point_re[120] = 'b1010010101111110;  // (-0.7071)
  assign point_re[121] = 'b1010100010000000;  // (-0.6836)
  assign point_re[122] = 'b1010101110011011;  // (-0.6593)
  assign point_re[123] = 'b1010111011001100;  // (-0.6344)
  assign point_re[124] = 'b1011001000010100;  // (-0.6088)
  assign point_re[125] = 'b1011010101110001;  // (-0.5825)
  assign point_re[126] = 'b1011100011100011;  // (-0.5556)
  assign point_re[127] = 'b1011110001101000;  // (-0.5281)
  assign point_re[128] = 'b1100000000000000;  // (-0.5000)
  assign point_re[129] = 'b1100001110101001;  // (-0.4714)
  assign point_re[130] = 'b1100011101100011;  // (-0.4423)
  assign point_re[131] = 'b1100101100101100;  // (-0.4127)
  assign point_re[132] = 'b1100111100000100;  // (-0.3827)
  assign point_re[133] = 'b1101001011101001;  // (-0.3523)
  assign point_re[134] = 'b1101011011011011;  // (-0.3214)
  assign point_re[135] = 'b1101101011011000;  // (-0.2903)
  assign point_re[136] = 'b1101111011011111;  // (-0.2588)
  assign point_re[137] = 'b1110001011101111;  // (-0.2271)
  assign point_re[138] = 'b1110011100000111;  // (-0.1951)
  assign point_re[139] = 'b1110101100100110;  // (-0.1629)
  assign point_re[140] = 'b1110111101001011;  // (-0.1305)
  assign point_re[141] = 'b1111001101110100;  // (-0.0980)
  assign point_re[142] = 'b1111011110100001;  // (-0.0654)
  assign point_re[143] = 'b1111101111010000;  // (-0.0327)
  assign point_re[144] = 'b0000000000000000;  // (-0.0000)
  assign point_re[145] = 'b0000010000110000;  // (0.0327)
  assign point_re[146] = 'b0000100001011111;  // (0.0654)
  assign point_re[147] = 'b0000110010001100;  // (0.0980)
  assign point_re[148] = 'b0001000010110101;  // (0.1305)
  assign point_re[149] = 'b0001010011011010;  // (0.1629)
  assign point_re[150] = 'b0001100011111001;  // (0.1951)
  assign point_re[151] = 'b0001110100010001;  // (0.2271)
  assign point_re[152] = 'b0010000100100001;  // (0.2588)
  assign point_re[153] = 'b0010010100101000;  // (0.2903)
  assign point_re[154] = 'b0010100100100101;  // (0.3214)
  assign point_re[155] = 'b0010110100010111;  // (0.3523)
  assign point_re[156] = 'b0011000011111100;  // (0.3827)
  assign point_re[157] = 'b0011010011010100;  // (0.4127)
  assign point_re[158] = 'b0011100010011101;  // (0.4423)
  assign point_re[159] = 'b0011110001010111;  // (0.4714)
  assign point_re[160] = 'b0100000000000000;  // (0.5000)
  assign point_re[161] = 'b0100001110011000;  // (0.5281)
  assign point_re[162] = 'b0100011100011101;  // (0.5556)
  assign point_re[163] = 'b0100101010001111;  // (0.5825)
  assign point_re[164] = 'b0100110111101100;  // (0.6088)
  assign point_re[165] = 'b0101000100110100;  // (0.6344)
  assign point_re[166] = 'b0101010001100101;  // (0.6593)
  assign point_re[167] = 'b0101011110000000;  // (0.6836)
  assign point_re[168] = 'b0101101010000010;  // (0.7071)
  assign point_re[169] = 'b0101110101101100;  // (0.7299)
  assign point_re[170] = 'b0110000000111100;  // (0.7518)
  assign point_re[171] = 'b0110001011110010;  // (0.7730)
  assign point_re[172] = 'b0110010110001101;  // (0.7934)
  assign point_re[173] = 'b0110100000001011;  // (0.8128)
  assign point_re[174] = 'b0110101001101110;  // (0.8315)
  assign point_re[175] = 'b0110110010110011;  // (0.8492)
  assign point_re[176] = 'b0110111011011010;  // (0.8660)
  assign point_re[177] = 'b0111000011100011;  // (0.8819)
  assign point_re[178] = 'b0111001011001101;  // (0.8969)
  assign point_re[179] = 'b0111010010010111;  // (0.9109)
  assign point_re[180] = 'b0111011001000010;  // (0.9239)
  assign point_re[181] = 'b0111011111001100;  // (0.9359)
  assign point_re[182] = 'b0111100100110101;  // (0.9469)
  assign point_re[183] = 'b0111101001111101;  // (0.9569)
  assign point_re[184] = 'b0111101110100011;  // (0.9659)
  assign point_re[185] = 'b0111110010101000;  // (0.9739)
  assign point_re[186] = 'b0111110110001010;  // (0.9808)
  assign point_re[187] = 'b0111111001001010;  // (0.9866)
  assign point_re[188] = 'b0111111011101000;  // (0.9914)
  assign point_re[189] = 'b0111111101100010;  // (0.9952)
  assign point_re[190] = 'b0111111110111010;  // (0.9979)
  assign point_re[191] = 'b0111111111101110;  // (0.9995)

  assign point_im[000] = 'b0000000000000000;  // (0.0000)
  assign point_im[001] = 'b0000010000110000;  // (0.0327)
  assign point_im[002] = 'b0000100001011111;  // (0.0654)
  assign point_im[003] = 'b0000110010001100;  // (0.0980)
  assign point_im[004] = 'b0001000010110101;  // (0.1305)
  assign point_im[005] = 'b0001010011011010;  // (0.1629)
  assign point_im[006] = 'b0001100011111001;  // (0.1951)
  assign point_im[007] = 'b0001110100010001;  // (0.2271)
  assign point_im[008] = 'b0010000100100001;  // (0.2588)
  assign point_im[009] = 'b0010010100101000;  // (0.2903)
  assign point_im[010] = 'b0010100100100101;  // (0.3214)
  assign point_im[011] = 'b0010110100010111;  // (0.3523)
  assign point_im[012] = 'b0011000011111100;  // (0.3827)
  assign point_im[013] = 'b0011010011010100;  // (0.4127)
  assign point_im[014] = 'b0011100010011101;  // (0.4423)
  assign point_im[015] = 'b0011110001010111;  // (0.4714)
  assign point_im[016] = 'b0100000000000000;  // (0.5000)
  assign point_im[017] = 'b0100001110011000;  // (0.5281)
  assign point_im[018] = 'b0100011100011101;  // (0.5556)
  assign point_im[019] = 'b0100101010001111;  // (0.5825)
  assign point_im[020] = 'b0100110111101100;  // (0.6088)
  assign point_im[021] = 'b0101000100110100;  // (0.6344)
  assign point_im[022] = 'b0101010001100101;  // (0.6593)
  assign point_im[023] = 'b0101011110000000;  // (0.6836)
  assign point_im[024] = 'b0101101010000010;  // (0.7071)
  assign point_im[025] = 'b0101110101101100;  // (0.7299)
  assign point_im[026] = 'b0110000000111100;  // (0.7518)
  assign point_im[027] = 'b0110001011110010;  // (0.7730)
  assign point_im[028] = 'b0110010110001101;  // (0.7934)
  assign point_im[029] = 'b0110100000001011;  // (0.8128)
  assign point_im[030] = 'b0110101001101110;  // (0.8315)
  assign point_im[031] = 'b0110110010110011;  // (0.8492)
  assign point_im[032] = 'b0110111011011010;  // (0.8660)
  assign point_im[033] = 'b0111000011100011;  // (0.8819)
  assign point_im[034] = 'b0111001011001101;  // (0.8969)
  assign point_im[035] = 'b0111010010010111;  // (0.9109)
  assign point_im[036] = 'b0111011001000010;  // (0.9239)
  assign point_im[037] = 'b0111011111001100;  // (0.9359)
  assign point_im[038] = 'b0111100100110101;  // (0.9469)
  assign point_im[039] = 'b0111101001111101;  // (0.9569)
  assign point_im[040] = 'b0111101110100011;  // (0.9659)
  assign point_im[041] = 'b0111110010101000;  // (0.9739)
  assign point_im[042] = 'b0111110110001010;  // (0.9808)
  assign point_im[043] = 'b0111111001001010;  // (0.9866)
  assign point_im[044] = 'b0111111011101000;  // (0.9914)
  assign point_im[045] = 'b0111111101100010;  // (0.9952)
  assign point_im[046] = 'b0111111110111010;  // (0.9979)
  assign point_im[047] = 'b0111111111101110;  // (0.9995)
  assign point_im[048] = 'b0111111111111111;  // (1.0000)
  assign point_im[049] = 'b0111111111101110;  // (0.9995)
  assign point_im[050] = 'b0111111110111010;  // (0.9979)
  assign point_im[051] = 'b0111111101100010;  // (0.9952)
  assign point_im[052] = 'b0111111011101000;  // (0.9914)
  assign point_im[053] = 'b0111111001001010;  // (0.9866)
  assign point_im[054] = 'b0111110110001010;  // (0.9808)
  assign point_im[055] = 'b0111110010101000;  // (0.9739)
  assign point_im[056] = 'b0111101110100011;  // (0.9659)
  assign point_im[057] = 'b0111101001111101;  // (0.9569)
  assign point_im[058] = 'b0111100100110101;  // (0.9469)
  assign point_im[059] = 'b0111011111001100;  // (0.9359)
  assign point_im[060] = 'b0111011001000010;  // (0.9239)
  assign point_im[061] = 'b0111010010010111;  // (0.9109)
  assign point_im[062] = 'b0111001011001101;  // (0.8969)
  assign point_im[063] = 'b0111000011100011;  // (0.8819)
  assign point_im[064] = 'b0110111011011010;  // (0.8660)
  assign point_im[065] = 'b0110110010110011;  // (0.8492)
  assign point_im[066] = 'b0110101001101110;  // (0.8315)
  assign point_im[067] = 'b0110100000001011;  // (0.8128)
  assign point_im[068] = 'b0110010110001101;  // (0.7934)
  assign point_im[069] = 'b0110001011110010;  // (0.7730)
  assign point_im[070] = 'b0110000000111100;  // (0.7518)
  assign point_im[071] = 'b0101110101101100;  // (0.7299)
  assign point_im[072] = 'b0101101010000010;  // (0.7071)
  assign point_im[073] = 'b0101011110000000;  // (0.6836)
  assign point_im[074] = 'b0101010001100101;  // (0.6593)
  assign point_im[075] = 'b0101000100110100;  // (0.6344)
  assign point_im[076] = 'b0100110111101100;  // (0.6088)
  assign point_im[077] = 'b0100101010001111;  // (0.5825)
  assign point_im[078] = 'b0100011100011101;  // (0.5556)
  assign point_im[079] = 'b0100001110011000;  // (0.5281)
  assign point_im[080] = 'b0100000000000000;  // (0.5000)
  assign point_im[081] = 'b0011110001010111;  // (0.4714)
  assign point_im[082] = 'b0011100010011101;  // (0.4423)
  assign point_im[083] = 'b0011010011010100;  // (0.4127)
  assign point_im[084] = 'b0011000011111100;  // (0.3827)
  assign point_im[085] = 'b0010110100010111;  // (0.3523)
  assign point_im[086] = 'b0010100100100101;  // (0.3214)
  assign point_im[087] = 'b0010010100101000;  // (0.2903)
  assign point_im[088] = 'b0010000100100001;  // (0.2588)
  assign point_im[089] = 'b0001110100010001;  // (0.2271)
  assign point_im[090] = 'b0001100011111001;  // (0.1951)
  assign point_im[091] = 'b0001010011011010;  // (0.1629)
  assign point_im[092] = 'b0001000010110101;  // (0.1305)
  assign point_im[093] = 'b0000110010001100;  // (0.0980)
  assign point_im[094] = 'b0000100001011111;  // (0.0654)
  assign point_im[095] = 'b0000010000110000;  // (0.0327)
  assign point_im[096] = 'b0000000000000000;  // (0.0000)
  assign point_im[097] = 'b1111101111010000;  // (-0.0327)
  assign point_im[098] = 'b1111011110100001;  // (-0.0654)
  assign point_im[099] = 'b1111001101110100;  // (-0.0980)
  assign point_im[100] = 'b1110111101001011;  // (-0.1305)
  assign point_im[101] = 'b1110101100100110;  // (-0.1629)
  assign point_im[102] = 'b1110011100000111;  // (-0.1951)
  assign point_im[103] = 'b1110001011101111;  // (-0.2271)
  assign point_im[104] = 'b1101111011011111;  // (-0.2588)
  assign point_im[105] = 'b1101101011011000;  // (-0.2903)
  assign point_im[106] = 'b1101011011011011;  // (-0.3214)
  assign point_im[107] = 'b1101001011101001;  // (-0.3523)
  assign point_im[108] = 'b1100111100000100;  // (-0.3827)
  assign point_im[109] = 'b1100101100101100;  // (-0.4127)
  assign point_im[110] = 'b1100011101100011;  // (-0.4423)
  assign point_im[111] = 'b1100001110101001;  // (-0.4714)
  assign point_im[112] = 'b1100000000000000;  // (-0.5000)
  assign point_im[113] = 'b1011110001101000;  // (-0.5281)
  assign point_im[114] = 'b1011100011100011;  // (-0.5556)
  assign point_im[115] = 'b1011010101110001;  // (-0.5825)
  assign point_im[116] = 'b1011001000010100;  // (-0.6088)
  assign point_im[117] = 'b1010111011001100;  // (-0.6344)
  assign point_im[118] = 'b1010101110011011;  // (-0.6593)
  assign point_im[119] = 'b1010100010000000;  // (-0.6836)
  assign point_im[120] = 'b1010010101111110;  // (-0.7071)
  assign point_im[121] = 'b1010001010010100;  // (-0.7299)
  assign point_im[122] = 'b1001111111000100;  // (-0.7518)
  assign point_im[123] = 'b1001110100001110;  // (-0.7730)
  assign point_im[124] = 'b1001101001110011;  // (-0.7934)
  assign point_im[125] = 'b1001011111110101;  // (-0.8128)
  assign point_im[126] = 'b1001010110010010;  // (-0.8315)
  assign point_im[127] = 'b1001001101001101;  // (-0.8492)
  assign point_im[128] = 'b1001000100100110;  // (-0.8660)
  assign point_im[129] = 'b1000111100011101;  // (-0.8819)
  assign point_im[130] = 'b1000110100110011;  // (-0.8969)
  assign point_im[131] = 'b1000101101101001;  // (-0.9109)
  assign point_im[132] = 'b1000100110111110;  // (-0.9239)
  assign point_im[133] = 'b1000100000110100;  // (-0.9359)
  assign point_im[134] = 'b1000011011001011;  // (-0.9469)
  assign point_im[135] = 'b1000010110000011;  // (-0.9569)
  assign point_im[136] = 'b1000010001011101;  // (-0.9659)
  assign point_im[137] = 'b1000001101011000;  // (-0.9739)
  assign point_im[138] = 'b1000001001110110;  // (-0.9808)
  assign point_im[139] = 'b1000000110110110;  // (-0.9866)
  assign point_im[140] = 'b1000000100011000;  // (-0.9914)
  assign point_im[141] = 'b1000000010011110;  // (-0.9952)
  assign point_im[142] = 'b1000000001000110;  // (-0.9979)
  assign point_im[143] = 'b1000000000010010;  // (-0.9995)
  assign point_im[144] = 'b1000000000000000;  // (-1.0000)
  assign point_im[145] = 'b1000000000010010;  // (-0.9995)
  assign point_im[146] = 'b1000000001000110;  // (-0.9979)
  assign point_im[147] = 'b1000000010011110;  // (-0.9952)
  assign point_im[148] = 'b1000000100011000;  // (-0.9914)
  assign point_im[149] = 'b1000000110110110;  // (-0.9866)
  assign point_im[150] = 'b1000001001110110;  // (-0.9808)
  assign point_im[151] = 'b1000001101011000;  // (-0.9739)
  assign point_im[152] = 'b1000010001011101;  // (-0.9659)
  assign point_im[153] = 'b1000010110000011;  // (-0.9569)
  assign point_im[154] = 'b1000011011001011;  // (-0.9469)
  assign point_im[155] = 'b1000100000110100;  // (-0.9359)
  assign point_im[156] = 'b1000100110111110;  // (-0.9239)
  assign point_im[157] = 'b1000101101101001;  // (-0.9109)
  assign point_im[158] = 'b1000110100110011;  // (-0.8969)
  assign point_im[159] = 'b1000111100011101;  // (-0.8819)
  assign point_im[160] = 'b1001000100100110;  // (-0.8660)
  assign point_im[161] = 'b1001001101001101;  // (-0.8492)
  assign point_im[162] = 'b1001010110010010;  // (-0.8315)
  assign point_im[163] = 'b1001011111110101;  // (-0.8128)
  assign point_im[164] = 'b1001101001110011;  // (-0.7934)
  assign point_im[165] = 'b1001110100001110;  // (-0.7730)
  assign point_im[166] = 'b1001111111000100;  // (-0.7518)
  assign point_im[167] = 'b1010001010010100;  // (-0.7299)
  assign point_im[168] = 'b1010010101111110;  // (-0.7071)
  assign point_im[169] = 'b1010100010000000;  // (-0.6836)
  assign point_im[170] = 'b1010101110011011;  // (-0.6593)
  assign point_im[171] = 'b1010111011001100;  // (-0.6344)
  assign point_im[172] = 'b1011001000010100;  // (-0.6088)
  assign point_im[173] = 'b1011010101110001;  // (-0.5825)
  assign point_im[174] = 'b1011100011100011;  // (-0.5556)
  assign point_im[175] = 'b1011110001101000;  // (-0.5281)
  assign point_im[176] = 'b1100000000000000;  // (-0.5000)
  assign point_im[177] = 'b1100001110101001;  // (-0.4714)
  assign point_im[178] = 'b1100011101100011;  // (-0.4423)
  assign point_im[179] = 'b1100101100101100;  // (-0.4127)
  assign point_im[180] = 'b1100111100000100;  // (-0.3827)
  assign point_im[181] = 'b1101001011101001;  // (-0.3523)
  assign point_im[182] = 'b1101011011011011;  // (-0.3214)
  assign point_im[183] = 'b1101101011011000;  // (-0.2903)
  assign point_im[184] = 'b1101111011011111;  // (-0.2588)
  assign point_im[185] = 'b1110001011101111;  // (-0.2271)
  assign point_im[186] = 'b1110011100000111;  // (-0.1951)
  assign point_im[187] = 'b1110101100100110;  // (-0.1629)
  assign point_im[188] = 'b1110111101001011;  // (-0.1305)
  assign point_im[189] = 'b1111001101110100;  // (-0.0980)
  assign point_im[190] = 'b1111011110100001;  // (-0.0654)
  assign point_im[191] = 'b1111101111010000;  // (-0.0327)

endmodule
