`timescale 1ns / 1ps

// `define TEST_F0
// `define TEST_F1
// `define TEST_F2
`define TEST_F3
// `define TEST_F4

/* PUCCH0
  PUCCH 0. [symStart nPUCCHSym] = [ 4  2]
  ack = 3 (2 bit), sr = 1 (1 bit)
  m0, nslot, nid = 5, 0, 512
  occi = 0
  mcs = 7

  PUCCH0 alpha * n + r = (10 *  0 + 15) mod 24 = 15/24 cyc. (-0.7071 + -0.7071i).   -0.7071 - 0.7071i
  PUCCH0 alpha * n + r = (10 *  1 +  9) mod 24 = 19/24 cyc. (00.2588 + -0.9659i).    0.2588 - 0.9659i
  PUCCH0 alpha * n + r = (10 *  2 +  9) mod 24 =  5/24 cyc. (00.2588 + 00.9659i).    0.2588 + 0.9659i
  PUCCH0 alpha * n + r = (10 *  3 +  3) mod 24 =  9/24 cyc. (-0.7071 + 00.7071i).   -0.7071 + 0.7071i
  PUCCH0 alpha * n + r = (10 *  4 + 15) mod 24 =  7/24 cyc. (-0.2588 + 00.9659i).   -0.2588 + 0.9659i
  PUCCH0 alpha * n + r = (10 *  5 +  9) mod 24 = 11/24 cyc. (-0.9659 + 00.2588i).   -0.9659 + 0.2588i
  PUCCH0 alpha * n + r = (10 *  6 + 21) mod 24 =  9/24 cyc. (-0.7071 + 00.7071i).   -0.7071 + 0.7071i
  PUCCH0 alpha * n + r = (10 *  7 +  3) mod 24 =  1/24 cyc. (00.9659 + 00.2588i).    0.9659 + 0.2588i
  PUCCH0 alpha * n + r = (10 *  8 +  9) mod 24 = 17/24 cyc. (-0.2588 + -0.9659i).   -0.2588 - 0.9659i
  PUCCH0 alpha * n + r = (10 *  9 + 15) mod 24 =  9/24 cyc. (-0.7071 + 00.7071i).   -0.7071 + 0.7071i
  PUCCH0 alpha * n + r = (10 * 10 +  9) mod 24 = 13/24 cyc. (-0.9659 + -0.2588i).   -0.9659 - 0.2588i
  PUCCH0 alpha * n + r = (10 * 11 + 15) mod 24 =  5/24 cyc. (00.2588 + 00.9659i).    0.2588 + 0.9659i
  PUCCH0 alpha * n + r = (10 *  0 + 15) mod 24 = 15/24 cyc. (-0.7071 + -0.7071i).   -0.7071 - 0.7071i
  PUCCH0 alpha * n + r = (10 *  1 +  9) mod 24 = 19/24 cyc. (00.2588 + -0.9659i).    0.2588 - 0.9659i
  PUCCH0 alpha * n + r = (10 *  2 +  9) mod 24 =  5/24 cyc. (00.2588 + 00.9659i).    0.2588 + 0.9659i
  PUCCH0 alpha * n + r = (10 *  3 +  3) mod 24 =  9/24 cyc. (-0.7071 + 00.7071i).   -0.7071 + 0.7071i
  PUCCH0 alpha * n + r = (10 *  4 + 15) mod 24 =  7/24 cyc. (-0.2588 + 00.9659i).   -0.2588 + 0.9659i
  PUCCH0 alpha * n + r = (10 *  5 +  9) mod 24 = 11/24 cyc. (-0.9659 + 00.2588i).   -0.9659 + 0.2588i
  PUCCH0 alpha * n + r = (10 *  6 + 21) mod 24 =  9/24 cyc. (-0.7071 + 00.7071i).   -0.7071 + 0.7071i
  PUCCH0 alpha * n + r = (10 *  7 +  3) mod 24 =  1/24 cyc. (00.9659 + 00.2588i).    0.9659 + 0.2588i
  PUCCH0 alpha * n + r = (10 *  8 +  9) mod 24 = 17/24 cyc. (-0.2588 + -0.9659i).   -0.2588 - 0.9659i
  PUCCH0 alpha * n + r = (10 *  9 + 15) mod 24 =  9/24 cyc. (-0.7071 + 00.7071i).   -0.7071 + 0.7071i
  PUCCH0 alpha * n + r = (10 * 10 +  9) mod 24 = 13/24 cyc. (-0.9659 + -0.2588i).   -0.9659 - 0.2588i
  PUCCH0 alpha * n + r = (10 * 11 + 15) mod 24 =  5/24 cyc. (00.2588 + 00.9659i).    0.2588 + 0.9659i
*/
/* PUCCH1
  |TESTBENCH  | y(n)  | wi(m)y(n) |

  PUCCH1 z = w + d + alpha * n + r = ( 0 + 15 + 14 *  0 + 15) mod 24 =  6/24 cyc. (00.0000 + 01.0000i). wi_phi =  0/24 cyc        -0.0000 + 1.0000i         -0.0000 + 1.0000i
  PUCCH1 z = w + d + alpha * n + r = ( 0 + 15 + 14 *  1 +  9) mod 24 = 14/24 cyc. (-0.8660 + -0.5000i). wi_phi =  0/24 cyc        -0.8660 - 0.5000i         -0.8660 - 0.5000i
  PUCCH1 z = w + d + alpha * n + r = ( 0 + 15 + 14 *  2 +  9) mod 24 =  4/24 cyc. (00.5000 + 00.8660i). wi_phi =  0/24 cyc         0.5000 + 0.8660i          0.5000 + 0.8660i
  PUCCH1 z = w + d + alpha * n + r = ( 0 + 15 + 14 *  3 +  3) mod 24 = 12/24 cyc. (-1.0000 + 00.0000i). wi_phi =  0/24 cyc        -1.0000 + 0.0000i         -1.0000 + 0.0000i
  PUCCH1 z = w + d + alpha * n + r = ( 0 + 15 + 14 *  4 + 15) mod 24 = 14/24 cyc. (-0.8660 + -0.5000i). wi_phi =  0/24 cyc        -0.8660 - 0.5000i         -0.8660 - 0.5000i
  PUCCH1 z = w + d + alpha * n + r = ( 0 + 15 + 14 *  5 +  9) mod 24 = 22/24 cyc. (00.8660 + -0.5000i). wi_phi =  0/24 cyc         0.8660 - 0.5000i          0.8660 - 0.5000i
  PUCCH1 z = w + d + alpha * n + r = ( 0 + 15 + 14 *  6 + 21) mod 24 =  0/24 cyc. (01.0000 + 00.0000i). wi_phi =  0/24 cyc         1.0000 - 0.0000i          1.0000 - 0.0000i
  PUCCH1 z = w + d + alpha * n + r = ( 0 + 15 + 14 *  7 +  3) mod 24 = 20/24 cyc. (00.5000 + -0.8660i). wi_phi =  0/24 cyc         0.5000 - 0.8660i          0.5000 - 0.8660i
  PUCCH1 z = w + d + alpha * n + r = ( 0 + 15 + 14 *  8 +  9) mod 24 = 16/24 cyc. (-0.5000 + -0.8660i). wi_phi =  0/24 cyc        -0.5000 - 0.8660i         -0.5000 - 0.8660i
  PUCCH1 z = w + d + alpha * n + r = ( 0 + 15 + 14 *  9 + 15) mod 24 = 12/24 cyc. (-1.0000 + 00.0000i). wi_phi =  0/24 cyc        -1.0000 - 0.0000i         -1.0000 - 0.0000i
  PUCCH1 z = w + d + alpha * n + r = ( 0 + 15 + 14 * 10 +  9) mod 24 = 20/24 cyc. (00.5000 + -0.8660i). wi_phi =  0/24 cyc         0.5000 - 0.8660i          0.5000 - 0.8660i
  PUCCH1 z = w + d + alpha * n + r = ( 0 + 15 + 14 * 11 + 15) mod 24 = 16/24 cyc. (-0.5000 + -0.8660i). wi_phi =  0/24 cyc        -0.5000 - 0.8660i         -0.5000 - 0.8660i
  PUCCH1 z = w + d + alpha * n + r = ( 8 + 15 + 22 *  0 + 15) mod 24 = 14/24 cyc. (-0.8660 + -0.5000i). wi_phi =  8/24 cyc        -0.0000 + 1.0000i         -0.8660 - 0.5000i
  PUCCH1 z = w + d + alpha * n + r = ( 8 + 15 + 22 *  1 +  9) mod 24 =  6/24 cyc. (00.0000 + 01.0000i). wi_phi =  8/24 cyc         0.8660 - 0.5000i          0.0000 + 1.0000i
  PUCCH1 z = w + d + alpha * n + r = ( 8 + 15 + 22 *  2 +  9) mod 24 =  4/24 cyc. (00.5000 + 00.8660i). wi_phi =  8/24 cyc         0.5000 - 0.8660i          0.5000 + 0.8660i
  PUCCH1 z = w + d + alpha * n + r = ( 8 + 15 + 22 *  3 +  3) mod 24 = 20/24 cyc. (00.5000 + -0.8660i). wi_phi =  8/24 cyc        -1.0000 + 0.0000i          0.5000 - 0.8660i
  PUCCH1 z = w + d + alpha * n + r = ( 8 + 15 + 22 *  4 + 15) mod 24 =  6/24 cyc. (00.0000 + 01.0000i). wi_phi =  8/24 cyc         0.8660 - 0.5000i          0.0000 + 1.0000i
  PUCCH1 z = w + d + alpha * n + r = ( 8 + 15 + 22 *  5 +  9) mod 24 = 22/24 cyc. (00.8660 + -0.5000i). wi_phi =  8/24 cyc        -0.8660 - 0.5000i          0.8660 - 0.5000i
  PUCCH1 z = w + d + alpha * n + r = ( 8 + 15 + 22 *  6 + 21) mod 24 =  8/24 cyc. (-0.5000 + 00.8660i). wi_phi =  8/24 cyc         1.0000 - 0.0000i         -0.5000 + 0.8660i
  PUCCH1 z = w + d + alpha * n + r = ( 8 + 15 + 22 *  7 +  3) mod 24 = 12/24 cyc. (-1.0000 + 00.0000i). wi_phi =  8/24 cyc         0.5000 + 0.8660i         -1.0000 + 0.0000i
  PUCCH1 z = w + d + alpha * n + r = ( 8 + 15 + 22 *  8 +  9) mod 24 = 16/24 cyc. (-0.5000 + -0.8660i). wi_phi =  8/24 cyc        -0.5000 + 0.8660i         -0.5000 - 0.8660i
  PUCCH1 z = w + d + alpha * n + r = ( 8 + 15 + 22 *  9 + 15) mod 24 = 20/24 cyc. (00.5000 + -0.8660i). wi_phi =  8/24 cyc        -1.0000 + 0.0000i          0.5000 - 0.8660i
  PUCCH1 z = w + d + alpha * n + r = ( 8 + 15 + 22 * 10 +  9) mod 24 = 12/24 cyc. (-1.0000 + 00.0000i). wi_phi =  8/24 cyc         0.5000 + 0.8660i         -1.0000 + 0.0000i
  PUCCH1 z = w + d + alpha * n + r = ( 8 + 15 + 22 * 11 + 15) mod 24 = 16/24 cyc. (-0.5000 + -0.8660i). wi_phi =  8/24 cyc        -0.5000 + 0.8660i         -0.5000 - 0.8660i
  PUCCH1 z = w + d + alpha * n + r = (16 + 15 + 20 *  0 + 15) mod 24 = 22/24 cyc. (00.8660 + -0.5000i). wi_phi = 16/24 cyc        -0.0000 + 1.0000i          0.8660 - 0.5000i
  PUCCH1 z = w + d + alpha * n + r = (16 + 15 + 20 *  1 +  9) mod 24 = 12/24 cyc. (-1.0000 + 00.0000i). wi_phi = 16/24 cyc         0.5000 - 0.8660i         -1.0000 + 0.0000i
  PUCCH1 z = w + d + alpha * n + r = (16 + 15 + 20 *  2 +  9) mod 24 =  8/24 cyc. (-0.5000 + 00.8660i). wi_phi = 16/24 cyc        -0.5000 - 0.8660i         -0.5000 + 0.8660i
  PUCCH1 z = w + d + alpha * n + r = (16 + 15 + 20 *  3 +  3) mod 24 = 22/24 cyc. (00.8660 + -0.5000i). wi_phi = 16/24 cyc         0.0000 + 1.0000i          0.8660 - 0.5000i
  PUCCH1 z = w + d + alpha * n + r = (16 + 15 + 20 *  4 + 15) mod 24 =  6/24 cyc. (00.0000 + 01.0000i). wi_phi = 16/24 cyc        -0.8660 - 0.5000i         -0.0000 + 1.0000i
  PUCCH1 z = w + d + alpha * n + r = (16 + 15 + 20 *  5 +  9) mod 24 = 20/24 cyc. (00.5000 + -0.8660i). wi_phi = 16/24 cyc         0.5000 + 0.8660i          0.5000 - 0.8660i
  PUCCH1 z = w + d + alpha * n + r = (16 + 15 + 20 *  6 + 21) mod 24 =  4/24 cyc. (00.5000 + 00.8660i). wi_phi = 16/24 cyc        -1.0000 + 0.0000i          0.5000 + 0.8660i
  PUCCH1 z = w + d + alpha * n + r = (16 + 15 + 20 *  7 +  3) mod 24 =  6/24 cyc. (00.0000 + 01.0000i). wi_phi = 16/24 cyc        -0.8660 - 0.5000i          0.0000 + 1.0000i
  PUCCH1 z = w + d + alpha * n + r = (16 + 15 + 20 *  8 +  9) mod 24 =  8/24 cyc. (-0.5000 + 00.8660i). wi_phi = 16/24 cyc        -0.5000 - 0.8660i         -0.5000 + 0.8660i
  PUCCH1 z = w + d + alpha * n + r = (16 + 15 + 20 *  9 + 15) mod 24 = 10/24 cyc. (-0.8660 + 00.5000i). wi_phi = 16/24 cyc         0.0000 - 1.0000i         -0.8660 + 0.5000i
  PUCCH1 z = w + d + alpha * n + r = (16 + 15 + 20 * 10 +  9) mod 24 =  0/24 cyc. (01.0000 + 00.0000i). wi_phi = 16/24 cyc        -0.5000 + 0.8660i          1.0000 + 0.0000i
  PUCCH1 z = w + d + alpha * n + r = (16 + 15 + 20 * 11 + 15) mod 24 =  2/24 cyc. (00.8660 + 00.5000i). wi_phi = 16/24 cyc        -0.8660 + 0.5000i          0.8660 + 0.5000i

  PUCCH 1. [symStart nPUCCHSym] = [ 4  7]
  ack = 1 (1 bit), sr = 0 (1 bit)
  m0, nslot, nid = 5, 3, 512
  occi = 1
  mcs = 0

  PUCCH1 z = w + d + alpha * n + r = ( 0 +  9 + 10 *  0 + 15) mod 24 =  0/24 cyc. (01.0000 + 00.0000i)          1.0000 + 0.0000i
  PUCCH1 z = w + d + alpha * n + r = ( 0 +  9 + 10 *  1 +  9) mod 24 =  4/24 cyc. (00.5000 + 00.8660i)          0.5000 + 0.8660i
  PUCCH1 z = w + d + alpha * n + r = ( 0 +  9 + 10 *  2 +  9) mod 24 = 14/24 cyc. (-0.8660 + -0.5000i)         -0.8660 - 0.5000i
  PUCCH1 z = w + d + alpha * n + r = ( 0 +  9 + 10 *  3 +  3) mod 24 = 18/24 cyc. (00.0000 + -1.0000i)         -0.0000 - 1.0000i
  PUCCH1 z = w + d + alpha * n + r = ( 0 +  9 + 10 *  4 + 15) mod 24 = 16/24 cyc. (-0.5000 + -0.8660i)         -0.5000 - 0.8660i
  PUCCH1 z = w + d + alpha * n + r = ( 0 +  9 + 10 *  5 +  9) mod 24 = 20/24 cyc. (00.5000 + -0.8660i)          0.5000 - 0.8660i
  PUCCH1 z = w + d + alpha * n + r = ( 0 +  9 + 10 *  6 + 21) mod 24 = 18/24 cyc. (00.0000 + -1.0000i)         -0.0000 - 1.0000i
  PUCCH1 z = w + d + alpha * n + r = ( 0 +  9 + 10 *  7 +  3) mod 24 = 10/24 cyc. (-0.8660 + 00.5000i)         -0.8660 + 0.5000i
  PUCCH1 z = w + d + alpha * n + r = ( 0 +  9 + 10 *  8 +  9) mod 24 =  2/24 cyc. (00.8660 + 00.5000i)          0.8660 + 0.5000i
  PUCCH1 z = w + d + alpha * n + r = ( 0 +  9 + 10 *  9 + 15) mod 24 = 18/24 cyc. (00.0000 + -1.0000i)          0.0000 - 1.0000i
  PUCCH1 z = w + d + alpha * n + r = ( 0 +  9 + 10 * 10 +  9) mod 24 = 22/24 cyc. (00.8660 + -0.5000i)          0.8660 - 0.5000i
  PUCCH1 z = w + d + alpha * n + r = ( 0 +  9 + 10 * 11 + 15) mod 24 = 14/24 cyc. (-0.8660 + -0.5000i)         -0.8660 - 0.5000i
  PUCCH1 z = w + d + alpha * n + r = (16 +  9 + 16 *  0 + 15) mod 24 = 16/24 cyc. (-0.5000 + -0.8660i)         -0.5000 - 0.8660i
  PUCCH1 z = w + d + alpha * n + r = (16 +  9 + 16 *  1 +  9) mod 24 =  2/24 cyc. (00.8660 + 00.5000i)          0.8660 + 0.5000i
  PUCCH1 z = w + d + alpha * n + r = (16 +  9 + 16 *  2 +  9) mod 24 = 18/24 cyc. (00.0000 + -1.0000i)         -0.0000 - 1.0000i
  PUCCH1 z = w + d + alpha * n + r = (16 +  9 + 16 *  3 +  3) mod 24 =  4/24 cyc. (00.5000 + 00.8660i)          0.5000 + 0.8660i
  PUCCH1 z = w + d + alpha * n + r = (16 +  9 + 16 *  4 + 15) mod 24 =  8/24 cyc. (-0.5000 + 00.8660i)         -0.5000 + 0.8660i
  PUCCH1 z = w + d + alpha * n + r = (16 +  9 + 16 *  5 +  9) mod 24 = 18/24 cyc. (00.0000 + -1.0000i)         -0.0000 - 1.0000i
  PUCCH1 z = w + d + alpha * n + r = (16 +  9 + 16 *  6 + 21) mod 24 = 22/24 cyc. (00.8660 + -0.5000i)          0.8660 - 0.5000i
  PUCCH1 z = w + d + alpha * n + r = (16 +  9 + 16 *  7 +  3) mod 24 = 20/24 cyc. (00.5000 + -0.8660i)          0.5000 - 0.8660i
  PUCCH1 z = w + d + alpha * n + r = (16 +  9 + 16 *  8 +  9) mod 24 = 18/24 cyc. (00.0000 + -1.0000i)         -0.0000 - 1.0000i
  PUCCH1 z = w + d + alpha * n + r = (16 +  9 + 16 *  9 + 15) mod 24 = 16/24 cyc. (-0.5000 + -0.8660i)         -0.5000 - 0.8660i
  PUCCH1 z = w + d + alpha * n + r = (16 +  9 + 16 * 10 +  9) mod 24 =  2/24 cyc. (00.8660 + 00.5000i)          0.8660 + 0.5000i
  PUCCH1 z = w + d + alpha * n + r = (16 +  9 + 16 * 11 + 15) mod 24 =  0/24 cyc. (01.0000 + 00.0000i)          1.0000 - 0.0000i
  PUCCH1 z = w + d + alpha * n + r = ( 8 +  9 +  6 *  0 + 15) mod 24 =  8/24 cyc. (-0.5000 + 00.8660i)         -0.5000 + 0.8660i
  PUCCH1 z = w + d + alpha * n + r = ( 8 +  9 +  6 *  1 +  9) mod 24 =  8/24 cyc. (-0.5000 + 00.8660i)         -0.5000 + 0.8660i
  PUCCH1 z = w + d + alpha * n + r = ( 8 +  9 +  6 *  2 +  9) mod 24 = 14/24 cyc. (-0.8660 + -0.5000i)         -0.8660 - 0.5000i
  PUCCH1 z = w + d + alpha * n + r = ( 8 +  9 +  6 *  3 +  3) mod 24 = 14/24 cyc. (-0.8660 + -0.5000i)         -0.8660 - 0.5000i
  PUCCH1 z = w + d + alpha * n + r = ( 8 +  9 +  6 *  4 + 15) mod 24 =  8/24 cyc. (-0.5000 + 00.8660i)         -0.5000 + 0.8660i
  PUCCH1 z = w + d + alpha * n + r = ( 8 +  9 +  6 *  5 +  9) mod 24 =  8/24 cyc. (-0.5000 + 00.8660i)         -0.5000 + 0.8660i
  PUCCH1 z = w + d + alpha * n + r = ( 8 +  9 +  6 *  6 + 21) mod 24 =  2/24 cyc. (00.8660 + 00.5000i)          0.8660 + 0.5000i
  PUCCH1 z = w + d + alpha * n + r = ( 8 +  9 +  6 *  7 +  3) mod 24 = 14/24 cyc. (-0.8660 + -0.5000i)         -0.8660 - 0.5000i
  PUCCH1 z = w + d + alpha * n + r = ( 8 +  9 +  6 *  8 +  9) mod 24 =  2/24 cyc. (00.8660 + 00.5000i)          0.8660 + 0.5000i
  PUCCH1 z = w + d + alpha * n + r = ( 8 +  9 +  6 *  9 + 15) mod 24 = 14/24 cyc. (-0.8660 + -0.5000i)         -0.8660 - 0.5000i
  PUCCH1 z = w + d + alpha * n + r = ( 8 +  9 +  6 * 10 +  9) mod 24 = 14/24 cyc. (-0.8660 + -0.5000i)         -0.8660 - 0.5000i
  PUCCH1 z = w + d + alpha * n + r = ( 8 +  9 +  6 * 11 + 15) mod 24 =  2/24 cyc. (00.8660 + 00.5000i)          0.8660 + 0.5000i

  PUCCH 1. [symStart nPUCCHSym] = [ 3  7]
  ack = 1 (2 bit), sr = 0 (1 bit)
  m0, nslot, nid = 5, 3, 512
  occi = 2
  mcs = 0
*/
/* PUCCH2
  PUCCH2 nid = 512, rnti = 56789 => cinit = 1860862464
  PUCCH2. d = QPSK(b( 0) ^ c( 0)) = QPSK(01) =  9/24 cyc (-0.7071 + 00.7071i)       -0.7071 + 0.7071i
  PUCCH2. d = QPSK(b( 1) ^ c( 1)) = QPSK(11) = 15/24 cyc (-0.7071 + -0.7071i)       -0.7071 - 0.7071i
  PUCCH2. d = QPSK(b( 2) ^ c( 2)) = QPSK(11) = 15/24 cyc (-0.7071 + -0.7071i)       -0.7071 - 0.7071i
  PUCCH2. d = QPSK(b( 3) ^ c( 3)) = QPSK(00) =  3/24 cyc (00.7071 + 00.7071i)        0.7071 + 0.7071i
  PUCCH2. d = QPSK(b( 4) ^ c( 4)) = QPSK(00) =  3/24 cyc (00.7071 + 00.7071i)        0.7071 + 0.7071i
  PUCCH2. d = QPSK(b( 5) ^ c( 5)) = QPSK(00) =  3/24 cyc (00.7071 + 00.7071i)        0.7071 + 0.7071i
  PUCCH2. d = QPSK(b( 6) ^ c( 6)) = QPSK(01) =  9/24 cyc (-0.7071 + 00.7071i)       -0.7071 + 0.7071i
  PUCCH2. d = QPSK(b( 7) ^ c( 7)) = QPSK(10) = 21/24 cyc (00.7071 + -0.7071i)        0.7071 - 0.7071i

  PUCCH2 nid = 512, rnti = 56789 => cinit = 1860862464
  sf, occi (n0), nIRB = 4, 2, 1 => n = (n0 + nIRB) mod sf = 3
  wn(i)d*d = w3(0)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i [ 0] d = QPSK(1) =  9/24 cyc
  wn(i)d*d = w3(1)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = w3(2)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = w3(3)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = w3(0)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i [ 1] d = QPSK(3) = 15/24 cyc
  wn(i)d*d = w3(1)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = w3(2)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = w3(3)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = w3(0)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i [ 2] d = QPSK(3) = 15/24 cyc
  wn(i)d*d = w3(1)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = w3(2)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = w3(3)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = w3(0)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i [ 3] d = QPSK(0) =  3/24 cyc
  wn(i)d*d = w3(1)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = w3(2)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = w3(3)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = w3(0)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i [ 4] d = QPSK(0) =  3/24 cyc
  wn(i)d*d = w3(1)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = w3(2)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = w3(3)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = w3(0)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i [ 5] d = QPSK(0) =  3/24 cyc
  wn(i)d*d = w3(1)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = w3(2)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = w3(3)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = w3(0)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i [ 6] d = QPSK(1) =  9/24 cyc
  wn(i)d*d = w3(1)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = w3(2)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = w3(3)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = w3(0)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i [ 7] d = QPSK(2) = 21/24 cyc
  wn(i)d*d = w3(1)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = w3(2)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = w3(3)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = w3(0)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i [ 8] d = QPSK(0) =  3/24 cyc
  wn(i)d*d = w3(1)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = w3(2)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = w3(3)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = w3(0)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i [ 9] d = QPSK(0) =  3/24 cyc
  wn(i)d*d = w3(1)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = w3(2)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = w3(3)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = w3(0)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i [10] d = QPSK(1) =  9/24 cyc
  wn(i)d*d = w3(1)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = w3(2)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = w3(3)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = w3(0)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i [11] d = QPSK(3) = 15/24 cyc
  wn(i)d*d = w3(1)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = w3(2)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = w3(3)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = w3(0)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i [12] d = QPSK(2) = 21/24 cyc
  wn(i)d*d = w3(1)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = w3(2)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = w3(3)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = w3(0)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i [13] d = QPSK(2) = 21/24 cyc
  wn(i)d*d = w3(1)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = w3(2)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = w3(3)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = w3(0)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i [14] d = QPSK(3) = 15/24 cyc
  wn(i)d*d = w3(1)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = w3(2)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = w3(3)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = w3(0)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i [15] d = QPSK(1) =  9/24 cyc
  wn(i)d*d = w3(1)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = w3(2)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = w3(3)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
*/

/* PUCCH3
  PUCCH3 nid = 512, rnti = 56789 => cinit = 1860862464
  Modulation = pi/2-BPSK. occi, sf = 2, 4. Mrb = 3

  Modulation symbols:
  [ 0] d = pi/2-BPSK(1) = 15/24 cyc
  [ 1] d = pi/2-BPSK(0) =  9/24 cyc
  [ 2] d = pi/2-BPSK(1) = 15/24 cyc
  [ 3] d = pi/2-BPSK(0) =  9/24 cyc
  [ 4] d = pi/2-BPSK(1) = 15/24 cyc
  [ 5] d = pi/2-BPSK(1) = 21/24 cyc
  [ 6] d = pi/2-BPSK(0) =  3/24 cyc
  [ 7] d = pi/2-BPSK(0) =  9/24 cyc
  [ 8] d = pi/2-BPSK(1) = 15/24 cyc
  [ 9] d = pi/2-BPSK(1) = 21/24 cyc
  [10] d = pi/2-BPSK(0) =  3/24 cyc
  [11] d = pi/2-BPSK(0) =  9/24 cyc
  [12] d = pi/2-BPSK(1) = 15/24 cyc
  [13] d = pi/2-BPSK(0) =  9/24 cyc
  [14] d = pi/2-BPSK(0) =  3/24 cyc
  [15] d = pi/2-BPSK(0) =  9/24 cyc
  [16] d = pi/2-BPSK(1) = 15/24 cyc
  [17] d = pi/2-BPSK(0) =  9/24 cyc
  [18] d = pi/2-BPSK(1) = 15/24 cyc
  [19] d = pi/2-BPSK(1) = 21/24 cyc
  [20] d = pi/2-BPSK(1) = 15/24 cyc
  [21] d = pi/2-BPSK(0) =  9/24 cyc
  [22] d = pi/2-BPSK(0) =  3/24 cyc
  [23] d = pi/2-BPSK(1) = 21/24 cyc
  [24] d = pi/2-BPSK(1) = 15/24 cyc
  [25] d = pi/2-BPSK(0) =  9/24 cyc
  [26] d = pi/2-BPSK(1) = 15/24 cyc
  [27] d = pi/2-BPSK(0) =  9/24 cyc
  [28] d = pi/2-BPSK(1) = 15/24 cyc
  [29] d = pi/2-BPSK(1) = 21/24 cyc
  [30] d = pi/2-BPSK(1) = 15/24 cyc
  [31] d = pi/2-BPSK(1) = 21/24 cyc
  [32] d = pi/2-BPSK(1) = 15/24 cyc
  [33] d = pi/2-BPSK(1) = 21/24 cyc
  [34] d = pi/2-BPSK(0) =  3/24 cyc
  [35] d = pi/2-BPSK(0) =  9/24 cyc
  [36] d = pi/2-BPSK(0) =  3/24 cyc
  [37] d = pi/2-BPSK(1) = 21/24 cyc
  [38] d = pi/2-BPSK(0) =  3/24 cyc
  [39] d = pi/2-BPSK(1) = 21/24 cyc
  [40] d = pi/2-BPSK(0) =  3/24 cyc
  [41] d = pi/2-BPSK(1) = 21/24 cyc
  [42] d = pi/2-BPSK(0) =  3/24 cyc
  [43] d = pi/2-BPSK(1) = 21/24 cyc
  [44] d = pi/2-BPSK(1) = 15/24 cyc
  [45] d = pi/2-BPSK(1) = 21/24 cyc
  [46] d = pi/2-BPSK(0) =  3/24 cyc
  [47] d = pi/2-BPSK(1) = 21/24 cyc
  [48] d = pi/2-BPSK(1) = 15/24 cyc
  [49] d = pi/2-BPSK(0) =  9/24 cyc
  [50] d = pi/2-BPSK(1) = 15/24 cyc
  [51] d = pi/2-BPSK(1) = 21/24 cyc
  [52] d = pi/2-BPSK(1) = 15/24 cyc
  [53] d = pi/2-BPSK(0) =  9/24 cyc
  [54] d = pi/2-BPSK(0) =  3/24 cyc
  [55] d = pi/2-BPSK(1) = 21/24 cyc
  [56] d = pi/2-BPSK(0) =  3/24 cyc
  [57] d = pi/2-BPSK(1) = 21/24 cyc
  [58] d = pi/2-BPSK(1) = 15/24 cyc
  [59] d = pi/2-BPSK(1) = 21/24 cyc
  [60] d = pi/2-BPSK(1) = 15/24 cyc
  [61] d = pi/2-BPSK(1) = 21/24 cyc
  [62] d = pi/2-BPSK(0) =  3/24 cyc
  [63] d = pi/2-BPSK(1) = 21/24 cyc
  [64] d = pi/2-BPSK(1) = 15/24 cyc
  [65] d = pi/2-BPSK(0) =  9/24 cyc
  [66] d = pi/2-BPSK(0) =  3/24 cyc
  [67] d = pi/2-BPSK(1) = 21/24 cyc
  [68] d = pi/2-BPSK(0) =  3/24 cyc
  [69] d = pi/2-BPSK(1) = 21/24 cyc
  [70] d = pi/2-BPSK(1) = 15/24 cyc
  [71] d = pi/2-BPSK(0) =  9/24 cyc

  wn(i)d*d = wx(0)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(1)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(1)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(1)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(1)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(1)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(1)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(1)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(1)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(1)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(1)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(1)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(1)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(1)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(1)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(1)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(1)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(1)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(1)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(1)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(1)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(1)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(1)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(1)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(1)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(1)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(1)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(1)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(1)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(1)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(1)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(1)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(1)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(1)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(1)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(1)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(1)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(1)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(1)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(1)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(1)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(1)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(1)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(1)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(1)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(1)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(1)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(1)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(1)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(1)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(1)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(1)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(1)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(1)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(1)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(1)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(1)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(1)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(1)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(1)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(1)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(1)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(1)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(1)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(1)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(1)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(1)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(1)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(1)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(1)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(1)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(1)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(1)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(2)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(2)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(2)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(2)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(2)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(2)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(2)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(2)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(2)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(2)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(2)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(2)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(2)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(2)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(2)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(2)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(2)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(2)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(2)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(2)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(2)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(2)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(2)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(2)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(2)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(2)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(2)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(2)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(2)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(2)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(2)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(2)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(2)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(2)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(2)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(2)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(2)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(2)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(2)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(2)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(2)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(2)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(2)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(2)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(2)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(2)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(2)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(2)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(2)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(2)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(2)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(2)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(2)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(2)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(2)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(2)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(2)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(2)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(2)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(2)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(2)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(2)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(2)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(2)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(2)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(2)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(2)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(2)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(2)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(2)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(2)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(2)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(3)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(3)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(3)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(3)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(3)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(3)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(3)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(3)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(3)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(3)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(3)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(3)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(3)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(3)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(3)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(3)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(3)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(3)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(3)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(3)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(3)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(3)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(3)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(3)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(3)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(3)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(3)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(3)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(3)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(3)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(3)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(3)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(3)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(3)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(3)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(3)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(3)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(3)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(3)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(3)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(3)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(3)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(3)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(3)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(3)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(3)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(3)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(3)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(3)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(3)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(3)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(3)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(3)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(3)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(3)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(3)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(3)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(3)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(3)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(3)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(3)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(3)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(3)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(3)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(3)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(3)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(3)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(3)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(3)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(3)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(3)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(3)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i


  PUCCH3 nid = 512, rnti = 56789 => cinit = 1860862464
  Modulation = pi/2-BPSK. occi, sf = 2, 0. Mrb = 3

  Modulation symbols:
  [ 0] d = pi/2-BPSK(1) = 15/24 cyc
  [ 1] d = pi/2-BPSK(0) =  9/24 cyc
  [ 2] d = pi/2-BPSK(1) = 15/24 cyc
  [ 3] d = pi/2-BPSK(0) =  9/24 cyc
  [ 4] d = pi/2-BPSK(1) = 15/24 cyc
  [ 5] d = pi/2-BPSK(1) = 21/24 cyc
  [ 6] d = pi/2-BPSK(0) =  3/24 cyc
  [ 7] d = pi/2-BPSK(0) =  9/24 cyc
  [ 8] d = pi/2-BPSK(1) = 15/24 cyc
  [ 9] d = pi/2-BPSK(1) = 21/24 cyc
  [10] d = pi/2-BPSK(0) =  3/24 cyc
  [11] d = pi/2-BPSK(0) =  9/24 cyc
  [12] d = pi/2-BPSK(1) = 15/24 cyc
  [13] d = pi/2-BPSK(0) =  9/24 cyc
  [14] d = pi/2-BPSK(0) =  3/24 cyc
  [15] d = pi/2-BPSK(0) =  9/24 cyc
  [16] d = pi/2-BPSK(1) = 15/24 cyc
  [17] d = pi/2-BPSK(0) =  9/24 cyc
  [18] d = pi/2-BPSK(1) = 15/24 cyc
  [19] d = pi/2-BPSK(1) = 21/24 cyc
  [20] d = pi/2-BPSK(1) = 15/24 cyc
  [21] d = pi/2-BPSK(0) =  9/24 cyc
  [22] d = pi/2-BPSK(0) =  3/24 cyc
  [23] d = pi/2-BPSK(1) = 21/24 cyc
  [24] d = pi/2-BPSK(1) = 15/24 cyc
  [25] d = pi/2-BPSK(0) =  9/24 cyc
  [26] d = pi/2-BPSK(1) = 15/24 cyc
  [27] d = pi/2-BPSK(0) =  9/24 cyc
  [28] d = pi/2-BPSK(1) = 15/24 cyc
  [29] d = pi/2-BPSK(1) = 21/24 cyc
  [30] d = pi/2-BPSK(1) = 15/24 cyc
  [31] d = pi/2-BPSK(1) = 21/24 cyc
  [32] d = pi/2-BPSK(1) = 15/24 cyc
  [33] d = pi/2-BPSK(1) = 21/24 cyc
  [34] d = pi/2-BPSK(0) =  3/24 cyc
  [35] d = pi/2-BPSK(0) =  9/24 cyc
  [36] d = pi/2-BPSK(0) =  3/24 cyc
  [37] d = pi/2-BPSK(1) = 21/24 cyc
  [38] d = pi/2-BPSK(0) =  3/24 cyc
  [39] d = pi/2-BPSK(1) = 21/24 cyc
  [40] d = pi/2-BPSK(0) =  3/24 cyc
  [41] d = pi/2-BPSK(1) = 21/24 cyc
  [42] d = pi/2-BPSK(0) =  3/24 cyc
  [43] d = pi/2-BPSK(1) = 21/24 cyc
  [44] d = pi/2-BPSK(1) = 15/24 cyc
  [45] d = pi/2-BPSK(1) = 21/24 cyc
  [46] d = pi/2-BPSK(0) =  3/24 cyc
  [47] d = pi/2-BPSK(1) = 21/24 cyc
  [48] d = pi/2-BPSK(1) = 15/24 cyc
  [49] d = pi/2-BPSK(0) =  9/24 cyc
  [50] d = pi/2-BPSK(1) = 15/24 cyc
  [51] d = pi/2-BPSK(1) = 21/24 cyc
  [52] d = pi/2-BPSK(1) = 15/24 cyc
  [53] d = pi/2-BPSK(0) =  9/24 cyc
  [54] d = pi/2-BPSK(0) =  3/24 cyc
  [55] d = pi/2-BPSK(1) = 21/24 cyc
  [56] d = pi/2-BPSK(0) =  3/24 cyc
  [57] d = pi/2-BPSK(1) = 21/24 cyc
  [58] d = pi/2-BPSK(1) = 15/24 cyc
  [59] d = pi/2-BPSK(1) = 21/24 cyc
  [60] d = pi/2-BPSK(1) = 15/24 cyc
  [61] d = pi/2-BPSK(1) = 21/24 cyc
  [62] d = pi/2-BPSK(0) =  3/24 cyc
  [63] d = pi/2-BPSK(1) = 21/24 cyc
  [64] d = pi/2-BPSK(1) = 15/24 cyc
  [65] d = pi/2-BPSK(0) =  9/24 cyc
  [66] d = pi/2-BPSK(0) =  3/24 cyc
  [67] d = pi/2-BPSK(1) = 21/24 cyc
  [68] d = pi/2-BPSK(0) =  3/24 cyc
  [69] d = pi/2-BPSK(1) = 21/24 cyc
  [70] d = pi/2-BPSK(1) = 15/24 cyc
  [71] d = pi/2-BPSK(0) =  9/24 cyc

  wn(i)d*d = wx(0)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d =  3/24 cyc (00.7071 + 00.7071)     0.7071 + 0.7071i
  wn(i)d*d = wx(0)*d = 21/24 cyc (00.7071 + -0.7071)     0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d = 15/24 cyc (-0.7071 + -0.7071)    -0.7071 - 0.7071i
  wn(i)d*d = wx(0)*d =  9/24 cyc (-0.7071 + 00.7071)    -0.7071 + 0.7071i
*/

// PUCCH 0 get nPUCCHSym(1-2) of alpha(s), starting from symStart(0-10)

module pucch_tb;

  // Parameters

  localparam nSlotSymb = 14;  //! (cyclic prefix (cp) == 'extended') ? 12 : 14
  localparam nRBSC = 12;

  localparam UNKNOWN = 16;

`ifdef TEST_F0
  /*
    PUCCH 0. [symStart nPUCCHSym] = [ 4  2]
    ack = 3 (2 bit), sr = 1 (1 bit)
    m0, nslot, nid = 5, 3, 512
    occi = 0
    mcs = 7
  */
  localparam VCD_FILE = "vcds/pucch0_tb.vcd";

  localparam test_pucch_format = 0;

  localparam test_symStart = 4;
  localparam test_nPUCCHSym = 2;  // nPUCCHSym = 7 => nSF = floor(nPUCCHSym/2) = 3

  localparam test_ack = 2'b11;  // ack = [bit1; bit0]
  localparam test_lenACK = 2;
  localparam test_sr = 1;
  localparam test_lenSR = 1;

  localparam test_m0 = 5;  // initialCS
  // localparam test_nslot = 3;
  localparam test_nslot = 0;
  localparam test_nid = 512;

  localparam lenUCI = 0;
`elsif TEST_F1
  /*
    PUCCH 1. [symStart nPUCCHSym] = [ 4  7]
    ack = 1 (1 bit), sr = 0 (1 bit)
    m0, nslot, nid = 5, 3, 512
    occi = 1
    mcs = 0
  */
  localparam VCD_FILE = "vcds/pucch1_tb.vcd";

  localparam test_pucch_format = 1;

  localparam test_symStart = 3;
  localparam test_nPUCCHSym = 7;  // nPUCCHSym = 7 => nSF = floor(nPUCCHSym/2) = 3

  localparam test_ack = 2'b01;  // ack = [bit1; bit0]
  localparam test_lenACK = 2;
  localparam test_sr = 0;
  localparam test_lenSR = 1;

  localparam test_m0 = 5;  // initialCS
  localparam test_nslot = 3;
  localparam test_nid = 512;

  localparam test_occi = 2;

  localparam lenUCI = 0;
`elsif TEST_F2
  localparam VCD_FILE = "vcds/pucch2_tb.vcd";
  localparam UCICW_FILE = "tb/pucch/uciCW_F2.txt";

  localparam test_pucch_format = 2;

  localparam test_rnti = 56789;  // F2
  localparam test_nid = 512;

  // n = (n0 + nIRB) mod sf
  localparam test_sf = 4;  // 2 or 4
  localparam test_occi = 2;  // n0
  localparam test_nIRB = 1;  // nIRB

  localparam lenUCI = 32;

  reg test_uciCW[0:lenUCI-1];
  integer test_uciCW_index;
  initial $readmemb(UCICW_FILE, test_uciCW);
`elsif TEST_F3
  localparam VCD_FILE = "vcds/pucch3_tb.vcd";
  localparam UCICW_FILE = "tb/pucch/uciCW_F3.txt";

  localparam test_pucch_format = 3;

  localparam test_rnti = 56789;  // F2
  localparam test_nid = 512;

  localparam test_sf = 0;  // 1 2 4
  localparam test_occi = 2;
  // localparam test_sf = 0;  // 1 2 4

  localparam test_Mrb = 3;  // F3
  localparam test_pi2bpsk_qpsk = 1;  // 1: pi/2 BPSK, 0: QPSK

  localparam lenUCI = 2 * (test_Mrb * nRBSC);

  reg test_uciCW[0:lenUCI-1];
  integer test_uciCW_index;
  initial $readmemb(UCICW_FILE, test_uciCW);
`elsif TEST_F4
  localparam VCD_FILE = "vcds/pucch4_tb.vcd";
  localparam UCICW_FILE = "tb/pucch/uciCW_F3.txt";

  localparam test_pucch_format = 4;

  localparam test_rnti = 56789;  // F2
  localparam test_nid = 512;

  localparam test_sf = 0;  // 1 2 4
  localparam test_occi = 2;
  // localparam test_sf = 0;  // 1 2 4

  localparam test_Mrb = 3;  // F3
  localparam test_pi2bpsk_qpsk = 1;  // 1: pi/2 BPSK, 0: QPSK

  localparam lenUCI = 2 * (test_Mrb * nRBSC);

  reg test_uciCW[0:lenUCI-1];
  integer test_uciCW_index;
  initial $readmemb(UCICW_FILE, test_uciCW);
`else

`endif

  initial begin
    begin
      $dumpfile(VCD_FILE);
      $dumpvars(10, pucch_dut);
      reset(3);
`ifdef TEST_F0
      test_f0f1(test_pucch_format,  //
                test_symStart, test_nPUCCHSym,  //
                test_ack, test_lenACK, test_sr, test_lenSR,  //
                test_m0, test_nslot, test_nid,  //
                0);
`elsif TEST_F1
      test_f0f1(test_pucch_format,  //
                test_symStart, test_nPUCCHSym,  //
                test_ack, test_lenACK, test_sr, test_lenSR,  //
                test_m0, test_nslot, test_nid,  //
                test_occi);
`elsif TEST_F2
      test_f2(test_pucch_format,  //
              test_nid, test_rnti,  //
              test_sf, test_occi, test_nIRB,  //
              lenUCI);
`elsif TEST_F3
      test_f234(test_pucch_format,  //
                test_nid, test_rnti,  //
                test_Mrb,  // No use
                lenUCI,  //
                test_pi2bpsk_qpsk,  //
                test_sf, test_occi);  //! The number of 2-bit value must be an integer multiple of (allocated number of subcarriers Msc = Mrb * nRBSC)
`elsif TEST_F4
      test_f234(test_pucch_format,  //
                test_nid, test_rnti,  //
                test_Mrb,  // No use
                lenUCI,  //
                test_pi2bpsk_qpsk,  //
                test_sf, test_occi);  //! The number of 2-bit value must be an integer multiple of (allocated number of subcarriers Msc = Mrb * nRBSC)
`else
`endif
      nop_clk(10);
      $finish;
    end
  end

  integer count_pucch = 0;
  string  disp_modulation;
  string  disp_output0;
  string  disp_output1;
  string  disp_output2;
  string  disp_output3;
  always @(posedge clk) begin
    if (o_valid) begin
      case (i_pucch_format)
        0: begin
          $write("PUCCH0 alpha * n + r = (%2d * %2d + %2d) mod 24 = %2d/24 cyc. (%07.4f + %07.4fi). ",  //
                 pucch_dut.alpha_cyc_24, pucch_dut.base_seq_n, pucch_dut.base_seq_cyc_24, pucch_dut.gen_parallel_pucch_234[0].point_cyc_24,  //
                 to_real(o_pucch_re[0]) / (2 ** 15), to_real(o_pucch_im[0]) / (2 ** 15));
          $display();
        end
        1: begin
          $write("PUCCH1 z = w + d + alpha * n + r = (%2d + %2d + %2d * %2d + %2d) mod 24 = %2d/24 cyc. (%07.4f + %07.4fi). ",  //
                 pucch_dut.spread_wi_phi_cyc_24, pucch_dut.cyc_24_modulation, pucch_dut.alpha_cyc_24, pucch_dut.base_seq_n, pucch_dut.base_seq_cyc_24, pucch_dut.gen_parallel_pucch_234[0].point_cyc_24,  //
                 to_real(o_pucch_re[0]) / (2 ** 15), to_real(o_pucch_im[0]) / (2 ** 15));
          // $display("wi_phi = %2d/24 cyc (is supported = %1b)", pucch_dut.spread_wi_phi_cyc_24, pucch_dut.spread_is_supported);
          $display();
        end
        2: begin
          count_pucch <= count_pucch + 1;
          $write("wn(i)d*d = w%1d(%1d)*d = %2d/24 cyc (%07.4f + %07.4f)",  //
                 (pucch_dut.i_occi + pucch_dut.i_nIRB) % pucch_dut.i_sf, 0, pucch_dut.gen_parallel_pucch_234[0].point_cyc_24,  //
                 to_real(pucch_dut.o_pucch_re[0]) / (2 ** 15), to_real(pucch_dut.o_pucch_im[0]) / (2 ** 15));
          $display(" [%2d] d = QPSK(%1d) = %2d/24 cyc",  //
                   count_pucch, pucch_dut.scrambler_scrambed_2bit, pucch_dut.d_qpsk);
          if (pucch_dut.gen_parallel_pucch_234[1].point_cyc_24) begin
            $display("wn(i)d*d = w%1d(%1d)*d = %2d/24 cyc (%07.4f + %07.4f)",  //
                     (pucch_dut.i_occi + pucch_dut.i_nIRB) % pucch_dut.i_sf, 1, pucch_dut.gen_parallel_pucch_234[1].point_cyc_24,  //
                     to_real(pucch_dut.o_pucch_re[1]) / (2 ** 15), to_real(pucch_dut.o_pucch_im[1]) / (2 ** 15));
          end
          if (pucch_dut.gen_parallel_pucch_234[2].point_cyc_24) begin
            $display("wn(i)d*d = w%1d(%1d)*d = %2d/24 cyc (%07.4f + %07.4f)",  //
                     (pucch_dut.i_occi + pucch_dut.i_nIRB) % pucch_dut.i_sf, 2, pucch_dut.gen_parallel_pucch_234[2].point_cyc_24,  //
                     to_real(pucch_dut.o_pucch_re[2]) / (2 ** 15), to_real(pucch_dut.o_pucch_im[2]) / (2 ** 15));
          end
          if (pucch_dut.gen_parallel_pucch_234[3].point_cyc_24) begin
            $display("wn(i)d*d = w%1d(%1d)*d = %2d/24 cyc (%07.4f + %07.4f)",  //
                     (pucch_dut.i_occi + pucch_dut.i_nIRB) % pucch_dut.i_sf, 3, pucch_dut.gen_parallel_pucch_234[3].point_cyc_24,  //
                     to_real(pucch_dut.o_pucch_re[3]) / (2 ** 15), to_real(pucch_dut.o_pucch_im[3]) / (2 ** 15));
          end
          // $display();
        end
        3, 4: begin
          count_pucch <= count_pucch + 1;
          $sformat(disp_modulation, "%s[%2d] d = %s(%1d) = %2d/24 cyc\n", disp_modulation,  //
                   count_pucch, pucch_dut.i_pi2bpsk_qpsk ? "pi/2-BPSK" : "QPSK", pucch_dut.i_pi2bpsk_qpsk ? pucch_dut.scrambler_scrambed_bit : pucch_dut.scrambler_scrambed_2bit, pucch_dut.i_pi2bpsk_qpsk ? pucch_dut.d_pi2bpsk : pucch_dut.d_qpsk);
          $sformat(disp_output0, "%swn(i)d*d = w%1d(%1d)*d = %2d/24 cyc (%07.4f + %07.4f)\n", disp_output0,  //
                   (pucch_dut.i_occi + pucch_dut.i_nIRB) % pucch_dut.i_sf, 0, pucch_dut.gen_parallel_pucch_234[0].point_cyc_24,  //
                   to_real(pucch_dut.o_pucch_re[0]) / (2 ** 15), to_real(pucch_dut.o_pucch_im[0]) / (2 ** 15));

          if (pucch_dut.gen_parallel_pucch_234[1].point_cyc_24) begin
            $sformat(disp_output1, "%swn(i)d*d = w%1d(%1d)*d = %2d/24 cyc (%07.4f + %07.4f)\n", disp_output1,  //
                     (pucch_dut.i_occi + pucch_dut.i_nIRB) % pucch_dut.i_sf, 1, pucch_dut.gen_parallel_pucch_234[1].point_cyc_24,  //
                     to_real(pucch_dut.o_pucch_re[1]) / (2 ** 15), to_real(pucch_dut.o_pucch_im[1]) / (2 ** 15));
          end
          if (pucch_dut.gen_parallel_pucch_234[2].point_cyc_24) begin
            $sformat(disp_output2, "%swn(i)d*d = w%1d(%1d)*d = %2d/24 cyc (%07.4f + %07.4f)\n", disp_output2,  //
                     (pucch_dut.i_occi + pucch_dut.i_nIRB) % pucch_dut.i_sf, 2, pucch_dut.gen_parallel_pucch_234[2].point_cyc_24,  //
                     to_real(pucch_dut.o_pucch_re[2]) / (2 ** 15), to_real(pucch_dut.o_pucch_im[2]) / (2 ** 15));
          end
          if (pucch_dut.gen_parallel_pucch_234[3].point_cyc_24) begin
            $sformat(disp_output3, "%swn(i)d*d = w%1d(%1d)*d = %2d/24 cyc (%07.4f + %07.4f)\n", disp_output3,  //
                     (pucch_dut.i_occi + pucch_dut.i_nIRB) % pucch_dut.i_sf, 3, pucch_dut.gen_parallel_pucch_234[3].point_cyc_24,  //
                     to_real(pucch_dut.o_pucch_re[3]) / (2 ** 15), to_real(pucch_dut.o_pucch_im[3]) / (2 ** 15));
          end
          if (count_pucch >= lenUCI - 1) begin
            $display("\nModulation symbols:\n%s", disp_modulation);
            $write("%s", disp_output0);
            $write("%s", disp_output1);
            $write("%s", disp_output2);
            $write("%s", disp_output3);
          end
        end
        default: begin
          $display("NOT A VALID PUCCH FORMAT (%1d)", pucch_dut.i_pucch_format);
        end
      endcase
    end
    if (o_done) begin
      nop_clk(10);
      $finish;
    end
  end

`ifdef TEST_F3
  task automatic test_f234;
    input integer pucch_format;
    input integer nid;
    input integer rnti;
    input integer Mrb;
    input integer get;
    input pi2bpsk_qpsk;
    input integer sf;
    input integer occi;
    integer uciCW;
    begin
      // @(negedge clk);
      i_pucch_format   = pucch_format;
      i_nid            = nid;
      i_rnti           = rnti;
      i_Mrb            = Mrb;
      i_pi2bpsk_qpsk   = pi2bpsk_qpsk;
      i_occi           = occi;
      i_sf             = sf;

      test_uciCW_index = 0;

      repeat (3) @(negedge clk);
      i_start = 1;
      @(negedge clk);
      i_start = 0;

      $display("PUCCH%1d nid = %1d, rnti = %1d => cinit = %1d", pucch_format, nid, rnti, pucch_dut.c_seq_gen_cinit);
      $display("Modulation = %s. occi, sf = %1d, %1d. Mrb = %1d", pi2bpsk_qpsk ? "pi/2-BPSK" : "QPSK", occi, sf, Mrb);

      repeat (get) begin
        i_uciCW = test_uciCW[test_uciCW_index];
        test_uciCW_index = test_uciCW_index + 1;

        i_uciCW_valid = 1;
        @(negedge clk);
        i_uciCW_valid = 0;
      end
    end
  endtask  //automatic
`endif

`ifdef TEST_F2
  task automatic test_f2;
    input integer pucch_format;
    input integer nid;
    input integer rnti;
    input integer sf;
    input integer occi;
    input integer nIRB;
    input integer get;
    integer uciCW;
    begin
      // @(negedge clk);
      i_pucch_format   = pucch_format;
      i_nid            = nid;
      i_rnti           = rnti;

      i_sf             = sf;
      i_occi           = occi;
      i_nIRB           = nIRB;

      test_uciCW_index = 0;

      repeat (3) @(negedge clk);
      i_start = 1;
      @(negedge clk);
      i_start = 0;

      $display("PUCCH2 nid = %1d, rnti = %1d => cinit = %1d", nid, rnti, pucch_dut.c_seq_gen_cinit);
      $display("sf, occi (n0), nIRB = %1d, %1d, %1d => n = (n0 + nIRB) mod sf = %1d", sf, occi, nIRB, (occi + nIRB) % sf);

      repeat (get) begin
        i_uciCW = test_uciCW[test_uciCW_index];
        test_uciCW_index = test_uciCW_index + 1;

        i_uciCW_valid = 1;
        @(negedge clk);
        i_uciCW_valid = 0;
      end
    end
  endtask  //automatic
`endif

  task automatic test_f0f1;
    input integer pucch_format;
    input integer symStart, nPUCCHSym;
    input integer ack, lenACK, sr, lenSR;
    input integer m0, nslot, nid;
    input integer occi;
    begin
      // @(negedge clk);
      i_pucch_format = pucch_format;
      i_symStart     = symStart;
      i_nPUCCHSym    = nPUCCHSym;
      i_ack          = ack;
      i_lenACK       = lenACK;
      i_sr           = sr;
      i_lenSR        = lenSR;
      i_m0           = m0;
      //   i_mcs          = mcs;
      i_nslot        = nslot;
      i_nid          = nid;
      i_occi         = occi;

      repeat (10) @(negedge clk);
      $display("PUCCH %1d. [symStart nPUCCHSym] = [%2d %2d]", pucch_format, symStart, nPUCCHSym);
      $display("ack = %1d (%1d bit), sr = %1d (%1d bit)", ack, lenACK, sr, lenSR);
      $display("m0, nslot, nid = %1d, %1d, %1d", m0, nslot, nid);
      $display("occi = %1d", occi);
      $display("mcs = %1d", pucch_dut.mcs);
      $display();

      i_start = 1;
      @(negedge clk);
      i_start = 0;

      @(negedge o_done);

    end
  endtask  //automatic

  // Ports
  reg                       clk = 0;
  reg                       rst = 0;
  reg         [        2:0] i_pucch_format;
  reg                       i_start = 0;
  reg         [        3:0] i_symStart;
  reg         [        3:0] i_nPUCCHSym;
  reg         [        1:0] i_ack;
  reg         [        1:0] i_lenACK;
  reg                       i_sr;
  reg                       i_lenSR;
  reg         [        3:0] i_m0;
  //   reg [3:0] i_mcs;
  reg         [        7:0] i_nslot;
  reg         [        9:0] i_nid;
  reg         [UNKNOWN-1:0] i_occi;

  reg         [       15:0] i_rnti;  //! [Format 2] Radio Network Temporary Identifier (0-65535)
  reg                       i_uciCW = 0;  //! [Format 2] Encoded UCI codeword as per TS 38.212 Section 6.3.1
  reg                       i_uciCW_valid = 0;  //! [Format 2] uciCW is valid and ready to continue generate PUCCH sequence
  reg         [        2:0] i_sf;
  reg         [UNKNOWN-1:0] i_nIRB;

  reg         [        4:0] i_Mrb;
  reg                       i_pi2bpsk_qpsk;

  wire signed [       15:0] o_pucch_re                                                                                     [0:3];
  wire signed [       15:0] o_pucch_im                                                                                     [0:3];
  wire                      o_valid;
  wire                      o_done;
  //

  pucch pucch_dut (
      .clk(clk),
      .rst(rst),

      .i_pucch_format(i_pucch_format),

      .i_start(i_start),

      .i_symStart (i_symStart),
      .i_nPUCCHSym(i_nPUCCHSym),

      .i_ack   (i_ack),
      .i_lenACK(i_lenACK),
      .i_sr    (i_sr),
      .i_lenSR (i_lenSR),

      .i_m0   (i_m0),
      //   .i_mcs  (i_mcs),
      .i_nslot(i_nslot),
      .i_nid  (i_nid),

      .i_occi(i_occi),

      .i_rnti       (i_rnti),
      .i_uciCW      (i_uciCW),
      .i_uciCW_valid(i_uciCW_valid),
      .i_sf         (i_sf),
      .i_nIRB       (i_nIRB),

      .i_Mrb(i_Mrb),
      .i_pi2bpsk_qpsk(i_pi2bpsk_qpsk),

      .o_pucch_re(o_pucch_re),
      .o_pucch_im(o_pucch_im),
      .o_valid   (o_valid),
      .o_done    (o_done)
  );

  task automatic reset;
    input integer clks;
    begin
      rst = 1;
      repeat (clks) @(negedge clk);
      rst = 0;
    end
  endtask  //automatic

  task automatic nop_clk;
    input integer clks;
    begin
      repeat (clks) @(posedge clk);
    end
  endtask  //automatic

  localparam CLK_PERIOD = 10;
  always #(CLK_PERIOD / 2) clk <= !clk;

  integer clk_count = 0;
  localparam MAX_CLK = 500;

  always @(posedge clk) begin
    clk_count <= clk_count + 1;
    if (clk_count > MAX_CLK) begin
      $display("MAX CLK");
      $finish;
    end
  end

  function real to_real;
    input signed [15:0] i_int;
    begin
      to_real = i_int;
    end
  endfunction

endmodule
